		when x"fe" => gain_n <= "000001000000111"; -- 80dB
		when x"fd" => gain_n <= "000001010001101"; -- 79dB
		when x"fc" => gain_n <= "000001100110111"; -- 78dB
		when x"fb" => gain_n <= "000010000001100"; -- 77dB
		when x"fa" => gain_n <= "000010100011000"; -- 76dB
		when x"f9" => gain_n <= "000011001101010"; -- 75dB
		when x"f8" => gain_n <= "000100000010011"; -- 74dB
		when x"f7" => gain_n <= "000101000101010"; -- 73dB
		when x"f6" => gain_n <= "000110011001100"; -- 72dB
		when x"f5" => gain_n <= "001000000011101"; -- 71dB
		when x"f4" => gain_n <= "001010001001001"; -- 70dB
		when x"f3" => gain_n <= "001100110001010"; -- 69dB
		when x"f2" => gain_n <= "010000000100110"; -- 68dB
		when x"f1" => gain_n <= "010100001111010"; -- 67dB
		when x"f0" => gain_n <= "010111010110111"; -- 66dB
		when x"ef" => gain_n <= "011001011101101"; -- 65dB
		when x"ee" => gain_n <= "011011100010100"; -- 64dB
		when x"ed" => gain_n <= "011101100101010"; -- 63dB
		when x"ec" => gain_n <= "011111100110000"; -- 62dB
		when x"eb" => gain_n <= "100001100100101"; -- 61dB
		when x"ea" => gain_n <= "100011100000111"; -- 60dB
		when x"e9" => gain_n <= "100101011010111"; -- 59dB
		when x"e8" => gain_n <= "100111010010100"; -- 58dB
		when x"e7" => gain_n <= "101001000111101"; -- 57dB
		when x"e6" => gain_n <= "101010111010001"; -- 56dB
		when x"e5" => gain_n <= "101100101001111"; -- 55dB
		when x"e4" => gain_n <= "101110010110111"; -- 54dB
		when x"e3" => gain_n <= "110000000000111"; -- 53dB
		when x"e2" => gain_n <= "110001100111111"; -- 52dB
		when x"e1" => gain_n <= "110011001011101"; -- 51dB
		when x"e0" => gain_n <= "110100101100001"; -- 50dB
		when x"df" => gain_n <= "110110001001001"; -- 49dB
		when x"de" => gain_n <= "110111100010100"; -- 48dB
		when x"dd" => gain_n <= "111000111000001"; -- 47dB
		when x"dc" => gain_n <= "111010001001111"; -- 46dB
		when x"db" => gain_n <= "111011010111011"; -- 45dB
		when x"da" => gain_n <= "111100100000100"; -- 44dB
		when x"d9" => gain_n <= "111101100101010"; -- 43dB
		when x"d8" => gain_n <= "111110100101001"; -- 42dB
		when x"d7" => gain_n <= "111111100000000"; -- 41dB
		when x"d6" => gain_n <= "111111111111111"; -- 40dB
		when x"d5" => gain_n <= "111111111111111"; -- 39dB
		when x"d4" => gain_n <= "111111111111111"; -- 38dB
		when x"d3" => gain_n <= "111111111111111"; -- 37dB
		when x"d2" => gain_n <= "111111111111111"; -- 36dB
		when x"d1" => gain_n <= "111111111111111"; -- 35dB
		when x"d0" => gain_n <= "111111111111111"; -- 34dB
		when x"cf" => gain_n <= "111111111111111"; -- 33dB
		when x"ce" => gain_n <= "111111111111111"; -- 32dB
		when x"cd" => gain_n <= "111111111111111"; -- 31dB
		when x"cc" => gain_n <= "111111111111111"; -- 30dB
		when x"cb" => gain_n <= "111111111111111"; -- 29dB
		when x"ca" => gain_n <= "111111111111111"; -- 28dB
		when x"c9" => gain_n <= "111111111111111"; -- 27dB
		when x"c8" => gain_n <= "111111111111111"; -- 26dB
		when x"c7" => gain_n <= "111111111111111"; -- 25dB
		when x"c6" => gain_n <= "111111111111111"; -- 24dB
		when x"c5" => gain_n <= "111111111111111"; -- 23dB
		when x"c4" => gain_n <= "111111111111111"; -- 22dB
		when x"c3" => gain_n <= "111111111111111"; -- 21dB
		when x"c2" => gain_n <= "111111111111111"; -- 20dB
		when x"c1" => gain_n <= "111111111111111"; -- 19dB
		when x"c0" => gain_n <= "111111111111111"; -- 18dB
		when x"bf" => gain_n <= "111111111111111"; -- 17dB
		when x"be" => gain_n <= "111111111111111"; -- 16dB
		when x"bd" => gain_n <= "111111111111111"; -- 15dB
		when x"bc" => gain_n <= "111111111111111"; -- 14dB
		when x"bb" => gain_n <= "111111111111111"; -- 13dB
		when x"ba" => gain_n <= "111111111111111"; -- 12dB
		when x"b9" => gain_n <= "111111111111111"; -- 11dB
		when x"b8" => gain_n <= "111111111111111"; -- 10dB
		when x"b7" => gain_n <= "111111111111111"; -- 9dB
		when x"b6" => gain_n <= "111111111111111"; -- 8dB
		when x"b5" => gain_n <= "111111111111111"; -- 7dB
		when x"b4" => gain_n <= "111111111111111"; -- 6dB
		when x"b3" => gain_n <= "111111111111111"; -- 5dB
		when x"b2" => gain_n <= "111111111111111"; -- 4dB
		when x"b1" => gain_n <= "111111111111111"; -- 3dB
		when x"b0" => gain_n <= "111111111111111"; -- 2dB
		when x"af" => gain_n <= "111111111111111"; -- 1dB
		when x"ae" => gain_n <= "111111111111111"; -- 0dB
