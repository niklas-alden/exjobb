        when x"08" => gain_n <= "000001000000111"; -- 90dB
        when x"07" => gain_n <= "000001010001101"; -- 89dB
        when x"06" => gain_n <= "000001100110111"; -- 88dB
        when x"05" => gain_n <= "000010000001100"; -- 87dB
        when x"04" => gain_n <= "000010100011000"; -- 86dB
        when x"03" => gain_n <= "000011001101010"; -- 85dB
        when x"02" => gain_n <= "000100000010011"; -- 84dB
        when x"01" => gain_n <= "000101000101010"; -- 83dB
        when x"00" => gain_n <= "000110011001100"; -- 82dB
        when x"ff" => gain_n <= "001000000011101"; -- 81dB
        when x"fe" => gain_n <= "001010001001001"; -- 80dB
        when x"fd" => gain_n <= "001101000011101"; -- 79dB
        when x"fc" => gain_n <= "001110100011100"; -- 78dB
        when x"fb" => gain_n <= "010000000010110"; -- 77dB
        when x"fa" => gain_n <= "010001100001101"; -- 76dB
        when x"f9" => gain_n <= "010010111111110"; -- 75dB
        when x"f8" => gain_n <= "010100011101011"; -- 74dB
        when x"f7" => gain_n <= "010101111010100"; -- 73dB
        when x"f6" => gain_n <= "010111010110111"; -- 72dB
        when x"f5" => gain_n <= "011000110010101"; -- 71dB
        when x"f4" => gain_n <= "011010001101110"; -- 70dB
        when x"f3" => gain_n <= "011011101000010"; -- 69dB
        when x"f2" => gain_n <= "011101000010000"; -- 68dB
        when x"f1" => gain_n <= "011110011010111"; -- 67dB
        when x"f0" => gain_n <= "011111110011001"; -- 66dB
        when x"ef" => gain_n <= "100001001010100"; -- 65dB
        when x"ee" => gain_n <= "100010100001000"; -- 64dB
        when x"ed" => gain_n <= "100011110110110"; -- 63dB
        when x"ec" => gain_n <= "100101001011100"; -- 62dB
        when x"eb" => gain_n <= "100110011111010"; -- 61dB
        when x"ea" => gain_n <= "100111110010001"; -- 60dB
        when x"e9" => gain_n <= "101001000100000"; -- 59dB
		when x"e8" => gain_n <= "101010010100101"; -- 58dB
        when x"e7" => gain_n <= "101011100100010"; -- 57dB
        when x"e6" => gain_n <= "101100110010110"; -- 56dB
        when x"e5" => gain_n <= "101101111111111"; -- 55dB
        when x"e4" => gain_n <= "101111001011110"; -- 54dB
        when x"e3" => gain_n <= "110000010110011"; -- 53dB
        when x"e2" => gain_n <= "110001011111100"; -- 52dB
        when x"e1" => gain_n <= "110010100111001"; -- 51dB
        when x"e0" => gain_n <= "110011101101010"; -- 50dB
        when x"df" => gain_n <= "110100110001110"; -- 49dB
        when x"de" => gain_n <= "110101110100100"; -- 48dB
        when x"dd" => gain_n <= "110110110101011"; -- 47dB
        when x"dc" => gain_n <= "110111110100100"; -- 46dB
        when x"db" => gain_n <= "111000110001100"; -- 45dB
        when x"da" => gain_n <= "111001101100011"; -- 44dB
        when x"d9" => gain_n <= "111010100101000"; -- 43dB
        when x"d8" => gain_n <= "111011011011010"; -- 42dB
        when x"d7" => gain_n <= "111100001111000"; -- 41dB
        when x"d6" => gain_n <= "111101000000001"; -- 40dB
        when x"d5" => gain_n <= "111101101110011"; -- 39dB
        when x"d4" => gain_n <= "111110011001101"; -- 38dB
        when x"d3" => gain_n <= "111111000001101"; -- 37dB
        when x"d2" => gain_n <= "111111100110011"; -- 36dB
        when x"d1" => gain_n <= "111111111111111"; -- 35dB
        when x"d0" => gain_n <= "111111111111111"; -- 34dB
        when x"cf" => gain_n <= "111111111111111"; -- 33dB
        when x"ce" => gain_n <= "111111111111111"; -- 32dB
        when x"cd" => gain_n <= "111111111111111"; -- 31dB
        when x"cc" => gain_n <= "111111111111111"; -- 30dB
        when x"cb" => gain_n <= "111111111111111"; -- 29dB
        when x"ca" => gain_n <= "111111111111111"; -- 28dB
        when x"c9" => gain_n <= "111111111111111"; -- 27dB
        when x"c8" => gain_n <= "111111111111111"; -- 26dB
        when x"c7" => gain_n <= "111111111111111"; -- 25dB
        when x"c6" => gain_n <= "111111111111111"; -- 24dB
        when x"c5" => gain_n <= "111111111111111"; -- 23dB
        when x"c4" => gain_n <= "111111111111111"; -- 22dB
        when x"c3" => gain_n <= "111111111111111"; -- 21dB
        when x"c2" => gain_n <= "111111111111111"; -- 20dB
        when x"c1" => gain_n <= "111111111111111"; -- 19dB
        when x"c0" => gain_n <= "111111111111111"; -- 18dB
        when x"bf" => gain_n <= "111111111111111"; -- 17dB
        when x"be" => gain_n <= "111111111111111"; -- 16dB
        when x"bd" => gain_n <= "111111111111111"; -- 15dB
        when x"bc" => gain_n <= "111111111111111"; -- 14dB
        when x"bb" => gain_n <= "111111111111111"; -- 13dB
        when x"ba" => gain_n <= "111111111111111"; -- 12dB
        when x"b9" => gain_n <= "111111111111111"; -- 11dB
        when x"b8" => gain_n <= "111111111111111"; -- 10dB
        when x"b7" => gain_n <= "111111111111111"; -- 9dB
        when x"b6" => gain_n <= "111111111111111"; -- 8dB
        when x"b5" => gain_n <= "111111111111111"; -- 7dB
        when x"b4" => gain_n <= "111111111111111"; -- 6dB
        when x"b3" => gain_n <= "111111111111111"; -- 5dB
        when x"b2" => gain_n <= "111111111111111"; -- 4dB
        when x"b1" => gain_n <= "111111111111111"; -- 3dB
        when x"b0" => gain_n <= "111111111111111"; -- 2dB
        when x"af" => gain_n <= "111111111111111"; -- 1dB
        when x"ae" => gain_n <= "111111111111111"; -- 0dB
        when x"ad" => gain_n <= "111111111111111"; -- -1dB
        when x"ac" => gain_n <= "111111111111111"; -- -2dB
        when x"ab" => gain_n <= "111111111111111"; -- -3dB
        when x"aa" => gain_n <= "111111111111111"; -- -4dB
        when x"a9" => gain_n <= "111111111111111"; -- -5dB
        when x"a8" => gain_n <= "111111111111111"; -- -6dB
        when x"a7" => gain_n <= "111111111111111"; -- -7dB
        when x"a6" => gain_n <= "111111111111111"; -- -8dB
        when x"a5" => gain_n <= "111111111111111"; -- -9dB
