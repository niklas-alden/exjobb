--------------------------------------------------------------------------------
-- Company: 
-- Engineer: Niklas Ald�n
--
-- Create Date:   17:00:43 03/25/2015
-- Design Name:   
-- Module Name:   D:/Google Drive/Exjobb/vhdl/agc_and_ac97/tb_top.vhd
-- Project Name:  agc_and_ac97
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: top
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
 
ENTITY tb_top IS
END tb_top;
 
ARCHITECTURE behavior OF tb_top IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT top
    PORT(
         clk : IN  std_logic;
         rstn : IN  std_logic;
         i_volume : IN  std_logic_vector(4 downto 0);
         i_SDATA_IN : IN  std_logic;
         o_SDATA_out : OUT  std_logic;
         o_SYNC : OUT  std_logic;
         o_RSTN : OUT  std_logic;
         i_BIT_CLK : IN  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal rstn : std_logic := '0';
   signal i_volume : std_logic_vector(4 downto 0) := (others => '0');
   signal i_SDATA_IN : std_logic := '0';
   signal i_BIT_CLK : std_logic := '0';

 	--Outputs
   signal o_SDATA_out : std_logic;
   signal o_SYNC : std_logic;
   signal o_RSTN : std_logic;

   -- Clock period definitions
   constant clk_period : time := 30.3 ns; -- 33MHz
   constant i_BIT_CLK_period : time := 81.38 ns; -- 12.288 MHz
   
   constant len : integer range 0 to 65535 := 20000;
   
	type t_sample is array(19 downto 0) of std_logic;
	type t_sample_matrix is array(0 to len-1) of t_sample;
	
	signal s : t_sample_matrix := (	
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"ffc00",-- -64
x"ffd00",-- -48
x"00000",-- 0
x"00200",-- 32
x"00100",-- 16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"00100",-- 16
x"00300",-- 48
x"00100",-- 16
x"fff00",-- -16
x"fff00",-- -16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffb00",-- -80
x"ffb00",-- -80
x"fff00",-- -16
x"00200",-- 32
x"00200",-- 32
x"ffe00",-- -32
x"ffc00",-- -64
x"fff00",-- -16
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"fff00",-- -16
x"00000",-- 0
x"00400",-- 64
x"00600",-- 96
x"00400",-- 64
x"00000",-- 0
x"ffd00",-- -48
x"ffe00",-- -32
x"00000",-- 0
x"00000",-- 0
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00200",-- 32
x"00200",-- 32
x"fff00",-- -16
x"ffd00",-- -48
x"00000",-- 0
x"00200",-- 32
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"ffc00",-- -64
x"ffc00",-- -64
x"fff00",-- -16
x"00200",-- 32
x"00100",-- 16
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"fff00",-- -16
x"00100",-- 16
x"00100",-- 16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffd00",-- -48
x"ffb00",-- -80
x"ffa00",-- -96
x"ffd00",-- -48
x"ffd00",-- -48
x"ffc00",-- -64
x"ffd00",-- -48
x"fff00",-- -16
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00300",-- 48
x"00500",-- 80
x"00300",-- 48
x"00000",-- 0
x"fff00",-- -16
x"00100",-- 16
x"00200",-- 32
x"00000",-- 0
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00200",-- 32
x"00100",-- 16
x"ffe00",-- -32
x"ffc00",-- -64
x"ffc00",-- -64
x"fff00",-- -16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"fff00",-- -16
x"00400",-- 64
x"00500",-- 80
x"00000",-- 0
x"ffc00",-- -64
x"ffc00",-- -64
x"fff00",-- -16
x"fff00",-- -16
x"ffd00",-- -48
x"ffc00",-- -64
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"ffd00",-- -48
x"ffd00",-- -48
x"00000",-- 0
x"00300",-- 48
x"00200",-- 32
x"fff00",-- -16
x"ffc00",-- -64
x"ffd00",-- -48
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00300",-- 48
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00400",-- 64
x"00500",-- 80
x"00300",-- 48
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00300",-- 48
x"00400",-- 64
x"00200",-- 32
x"fff00",-- -16
x"ffc00",-- -64
x"ffc00",-- -64
x"ffe00",-- -32
x"00000",-- 0
x"00200",-- 32
x"00300",-- 48
x"00000",-- 0
x"ffe00",-- -32
x"ffe00",-- -32
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"ffe00",-- -32
x"ffd00",-- -48
x"fff00",-- -16
x"00200",-- 32
x"00500",-- 80
x"00300",-- 48
x"00100",-- 16
x"00000",-- 0
x"00200",-- 32
x"00500",-- 80
x"00300",-- 48
x"00000",-- 0
x"ffe00",-- -32
x"00100",-- 16
x"00400",-- 64
x"00200",-- 32
x"ffe00",-- -32
x"fff00",-- -16
x"00200",-- 32
x"00400",-- 64
x"00300",-- 48
x"00300",-- 48
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00500",-- 80
x"00600",-- 96
x"00300",-- 48
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00200",-- 32
x"00100",-- 16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"ffe00",-- -32
x"ffd00",-- -48
x"fff00",-- -16
x"00200",-- 32
x"00300",-- 48
x"00100",-- 16
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"00100",-- 16
x"00300",-- 48
x"00000",-- 0
x"ffc00",-- -64
x"ffe00",-- -32
x"00300",-- 48
x"00400",-- 64
x"00200",-- 32
x"00000",-- 0
x"00000",-- 0
x"00200",-- 32
x"00400",-- 64
x"00400",-- 64
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00300",-- 48
x"00200",-- 32
x"00000",-- 0
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00200",-- 32
x"00300",-- 48
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00100",-- 16
x"00100",-- 16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"ffd00",-- -48
x"fff00",-- -16
x"00200",-- 32
x"00100",-- 16
x"ffe00",-- -32
x"ffe00",-- -32
x"00200",-- 32
x"00600",-- 96
x"00400",-- 64
x"fff00",-- -16
x"ffc00",-- -64
x"ffe00",-- -32
x"00200",-- 32
x"00200",-- 32
x"fff00",-- -16
x"ffd00",-- -48
x"ffe00",-- -32
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"ffd00",-- -48
x"ffd00",-- -48
x"fff00",-- -16
x"fff00",-- -16
x"ffc00",-- -64
x"ffa00",-- -96
x"ffc00",-- -64
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"ffd00",-- -48
x"ffd00",-- -48
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00200",-- 32
x"00100",-- 16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00200",-- 32
x"00300",-- 48
x"00100",-- 16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00200",-- 32
x"00200",-- 32
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00200",-- 32
x"00300",-- 48
x"00000",-- 0
x"ffd00",-- -48
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00200",-- 32
x"00400",-- 64
x"00400",-- 64
x"00300",-- 48
x"00100",-- 16
x"ffe00",-- -32
x"ffd00",-- -48
x"fff00",-- -16
x"00200",-- 32
x"00300",-- 48
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00300",-- 48
x"00300",-- 48
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00300",-- 48
x"00400",-- 64
x"00300",-- 48
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00300",-- 48
x"00200",-- 32
x"fff00",-- -16
x"ffd00",-- -48
x"ffd00",-- -48
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00100",-- 16
x"00300",-- 48
x"00400",-- 64
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00100",-- 16
x"00300",-- 48
x"00300",-- 48
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00300",-- 48
x"00300",-- 48
x"00000",-- 0
x"ffd00",-- -48
x"ffe00",-- -32
x"00100",-- 16
x"00200",-- 32
x"00000",-- 0
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"ffc00",-- -64
x"ffc00",-- -64
x"fff00",-- -16
x"00100",-- 16
x"00000",-- 0
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffc00",-- -64
x"ffd00",-- -48
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"ffd00",-- -48
x"ffd00",-- -48
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"ffc00",-- -64
x"ffd00",-- -48
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffd00",-- -48
x"fff00",-- -16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"fff00",-- -16
x"00200",-- 32
x"00300",-- 48
x"00300",-- 48
x"00200",-- 32
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00300",-- 48
x"00400",-- 64
x"00200",-- 32
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00400",-- 64
x"00400",-- 64
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00200",-- 32
x"00400",-- 64
x"00300",-- 48
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00200",-- 32
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"ffe00",-- -32
x"ffc00",-- -64
x"fff00",-- -16
x"00200",-- 32
x"00200",-- 32
x"fff00",-- -16
x"ffc00",-- -64
x"ffd00",-- -48
x"00000",-- 0
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"fff00",-- -16
x"00200",-- 32
x"00300",-- 48
x"00100",-- 16
x"fff00",-- -16
x"fff00",-- -16
x"00100",-- 16
x"00300",-- 48
x"00300",-- 48
x"00000",-- 0
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00100",-- 16
x"00000",-- 0
x"ffd00",-- -48
x"ffc00",-- -64
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00300",-- 48
x"00100",-- 16
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"ffd00",-- -48
x"ffb00",-- -80
x"ffc00",-- -64
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffb00",-- -80
x"ffb00",-- -80
x"ffd00",-- -48
x"ffd00",-- -48
x"ffc00",-- -64
x"ffb00",-- -80
x"ffa00",-- -96
x"ffb00",-- -80
x"ffd00",-- -48
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"fff00",-- -16
x"ffd00",-- -48
x"ffe00",-- -32
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00300",-- 48
x"00100",-- 16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"00100",-- 16
x"00300",-- 48
x"00100",-- 16
x"ffe00",-- -32
x"ffc00",-- -64
x"fff00",-- -16
x"00100",-- 16
x"00100",-- 16
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00200",-- 32
x"00100",-- 16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00300",-- 48
x"00400",-- 64
x"00500",-- 80
x"00400",-- 64
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00300",-- 48
x"00200",-- 32
x"00000",-- 0
x"00100",-- 16
x"00300",-- 48
x"00300",-- 48
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00200",-- 32
x"00400",-- 64
x"00100",-- 16
x"ffe00",-- -32
x"fff00",-- -16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffd00",-- -48
x"ffc00",-- -64
x"ffc00",-- -64
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00200",-- 32
x"00400",-- 64
x"00300",-- 48
x"00200",-- 32
x"00200",-- 32
x"00400",-- 64
x"00500",-- 80
x"00400",-- 64
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"fff00",-- -16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"ffe00",-- -32
x"fff00",-- -16
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"00100",-- 16
x"00200",-- 32
x"00000",-- 0
x"ffd00",-- -48
x"ffd00",-- -48
x"fff00",-- -16
x"00100",-- 16
x"00100",-- 16
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"00000",-- 0
x"00300",-- 48
x"00300",-- 48
x"00200",-- 32
x"00000",-- 0
x"fff00",-- -16
x"00100",-- 16
x"00300",-- 48
x"00200",-- 32
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"fff00",-- -16
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00000",-- 0
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"fff00",-- -16
x"ffc00",-- -64
x"ffb00",-- -80
x"ffe00",-- -32
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"ffd00",-- -48
x"ffb00",-- -80
x"ffc00",-- -64
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffc00",-- -64
x"ffc00",-- -64
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffc00",-- -64
x"ffb00",-- -80
x"ffd00",-- -48
x"fff00",-- -16
x"fff00",-- -16
x"ffc00",-- -64
x"ffa00",-- -96
x"ffc00",-- -64
x"00000",-- 0
x"00100",-- 16
x"fff00",-- -16
x"ffc00",-- -64
x"ffc00",-- -64
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"fff00",-- -16
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffc00",-- -64
x"ffc00",-- -64
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffb00",-- -80
x"ffc00",-- -64
x"fff00",-- -16
x"fff00",-- -16
x"ffc00",-- -64
x"ffc00",-- -64
x"00000",-- 0
x"00200",-- 32
x"00100",-- 16
x"ffe00",-- -32
x"ffc00",-- -64
x"ffd00",-- -48
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"fff00",-- -16
x"ffe00",-- -32
x"00100",-- 16
x"00300",-- 48
x"00200",-- 32
x"ffe00",-- -32
x"ffd00",-- -48
x"fff00",-- -16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00300",-- 48
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00300",-- 48
x"00300",-- 48
x"00300",-- 48
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00200",-- 32
x"00400",-- 64
x"00400",-- 64
x"00200",-- 32
x"00000",-- 0
x"00100",-- 16
x"00300",-- 48
x"00500",-- 80
x"00200",-- 32
x"fff00",-- -16
x"ffd00",-- -48
x"fff00",-- -16
x"00200",-- 32
x"00100",-- 16
x"ffe00",-- -32
x"ffc00",-- -64
x"ffb00",-- -80
x"ffe00",-- -32
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"ffc00",-- -64
x"ffd00",-- -48
x"ffe00",-- -32
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"fff00",-- -16
x"ffd00",-- -48
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"ffd00",-- -48
x"ffd00",-- -48
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00300",-- 48
x"00200",-- 32
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00100",-- 16
x"00100",-- 16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"ffd00",-- -48
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"ffd00",-- -48
x"ffc00",-- -64
x"ffc00",-- -64
x"ffc00",-- -64
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffc00",-- -64
x"ffc00",-- -64
x"ffc00",-- -64
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"fff00",-- -16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffb00",-- -80
x"ffb00",-- -80
x"ffc00",-- -64
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00100",-- 16
x"00200",-- 32
x"00300",-- 48
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00300",-- 48
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"fff00",-- -16
x"00200",-- 32
x"00300",-- 48
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"ffd00",-- -48
x"ffe00",-- -32
x"00000",-- 0
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00300",-- 48
x"00300",-- 48
x"00200",-- 32
x"00200",-- 32
x"00300",-- 48
x"00300",-- 48
x"00300",-- 48
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00300",-- 48
x"00100",-- 16
x"fff00",-- -16
x"fff00",-- -16
x"00100",-- 16
x"00300",-- 48
x"00100",-- 16
x"fff00",-- -16
x"fff00",-- -16
x"00100",-- 16
x"00300",-- 48
x"00300",-- 48
x"00000",-- 0
x"ffe00",-- -32
x"fff00",-- -16
x"00100",-- 16
x"00200",-- 32
x"00000",-- 0
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"ffd00",-- -48
x"ffd00",-- -48
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"fff00",-- -16
x"ffd00",-- -48
x"ffd00",-- -48
x"fff00",-- -16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"ffd00",-- -48
x"ffc00",-- -64
x"ffd00",-- -48
x"fff00",-- -16
x"00000",-- 0
x"ffe00",-- -32
x"ffc00",-- -64
x"ffc00",-- -64
x"fff00",-- -16
x"00100",-- 16
x"00100",-- 16
x"ffe00",-- -32
x"ffc00",-- -64
x"ffd00",-- -48
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"ffd00",-- -48
x"ffc00",-- -64
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"00100",-- 16
x"00200",-- 32
x"00000",-- 0
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"fff00",-- -16
x"ffd00",-- -48
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"fff00",-- -16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"fff00",-- -16
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffc00",-- -64
x"ffe00",-- -32
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffc00",-- -64
x"ffc00",-- -64
x"ffd00",-- -48
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"fff00",-- -16
x"ffc00",-- -64
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffc00",-- -64
x"ffd00",-- -48
x"ffd00",-- -48
x"ffc00",-- -64
x"ffc00",-- -64
x"ffc00",-- -64
x"ffd00",-- -48
x"ffc00",-- -64
x"ffc00",-- -64
x"ffc00",-- -64
x"ffc00",-- -64
x"ffc00",-- -64
x"ffd00",-- -48
x"ffd00",-- -48
x"ffc00",-- -64
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffc00",-- -64
x"ffc00",-- -64
x"ffb00",-- -80
x"ffa00",-- -96
x"ffa00",-- -96
x"ff900",-- -112
x"ff900",-- -112
x"ff900",-- -112
x"ff800",-- -128
x"ff800",-- -128
x"ff800",-- -128
x"ff900",-- -112
x"ff800",-- -128
x"ff900",-- -112
x"ff900",-- -112
x"ffa00",-- -96
x"ffa00",-- -96
x"ffc00",-- -64
x"ffc00",-- -64
x"ffd00",-- -48
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00300",-- 48
x"00400",-- 64
x"00500",-- 80
x"00500",-- 80
x"00700",-- 112
x"00700",-- 112
x"00800",-- 128
x"00900",-- 144
x"00900",-- 144
x"00900",-- 144
x"00a00",-- 160
x"00b00",-- 176
x"00b00",-- 176
x"00b00",-- 176
x"00b00",-- 176
x"00a00",-- 160
x"00800",-- 128
x"00500",-- 80
x"00200",-- 32
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffd00",-- -48
x"ff800",-- -128
x"ff400",-- -192
x"ff200",-- -224
x"ff100",-- -240
x"ff000",-- -256
x"fed00",-- -304
x"fea00",-- -352
x"fe700",-- -400
x"fe700",-- -400
x"fe900",-- -368
x"fea00",-- -352
x"fea00",-- -352
x"fe900",-- -368
x"fea00",-- -352
x"fed00",-- -304
x"ff100",-- -240
x"ff500",-- -176
x"ff800",-- -128
x"ffb00",-- -80
x"ffe00",-- -32
x"00200",-- 32
x"00500",-- 80
x"00900",-- 144
x"00d00",-- 208
x"01000",-- 256
x"01200",-- 288
x"01400",-- 320
x"01600",-- 352
x"01900",-- 400
x"01c00",-- 448
x"01e00",-- 480
x"01e00",-- 480
x"01e00",-- 480
x"01f00",-- 496
x"02000",-- 512
x"02000",-- 512
x"02000",-- 512
x"01600",-- 352
x"00200",-- 32
x"ffc00",-- -64
x"00800",-- 128
x"01200",-- 288
x"00600",-- 96
x"ff200",-- -224
x"fe500",-- -432
x"fe100",-- -496
x"fe800",-- -384
x"ff200",-- -224
x"feb00",-- -336
x"fd600",-- -672
x"fce00",-- -800
x"fd700",-- -656
x"fe100",-- -496
x"fe500",-- -432
x"fe900",-- -368
x"fe700",-- -400
x"fe300",-- -464
x"feb00",-- -336
x"ffc00",-- -64
x"00400",-- 64
x"00900",-- 144
x"01100",-- 272
x"01400",-- 320
x"01200",-- 288
x"01600",-- 352
x"02000",-- 512
x"02400",-- 576
x"02600",-- 608
x"02500",-- 592
x"01c00",-- 448
x"01300",-- 304
x"01400",-- 320
x"01800",-- 384
x"01400",-- 320
x"00a00",-- 160
x"fff00",-- -16
x"ff400",-- -192
x"fee00",-- -288
x"ff000",-- -256
x"fef00",-- -272
x"fe700",-- -400
x"fde00",-- -544
x"fd900",-- -624
x"fd700",-- -656
x"fd900",-- -624
x"fdf00",-- -528
x"fe200",-- -480
x"fe200",-- -480
x"fe200",-- -480
x"fe500",-- -432
x"feb00",-- -336
x"ff300",-- -208
x"ffd00",-- -48
x"00300",-- 48
x"00400",-- 64
x"00600",-- 96
x"00c00",-- 192
x"01200",-- 288
x"01900",-- 400
x"01d00",-- 464
x"01d00",-- 464
x"01a00",-- 416
x"01800",-- 384
x"01900",-- 400
x"01b00",-- 432
x"01a00",-- 416
x"01600",-- 352
x"00f00",-- 240
x"00900",-- 144
x"00500",-- 80
x"00300",-- 48
x"00000",-- 0
x"ffc00",-- -64
x"ff700",-- -144
x"ff100",-- -240
x"fed00",-- -304
x"fec00",-- -320
x"fec00",-- -320
x"fed00",-- -304
x"fec00",-- -320
x"feb00",-- -336
x"feb00",-- -336
x"fec00",-- -320
x"ff000",-- -256
x"ff500",-- -176
x"ff900",-- -112
x"ffc00",-- -64
x"ffd00",-- -48
x"fff00",-- -16
x"00300",-- 48
x"00900",-- 144
x"00d00",-- 208
x"00f00",-- 240
x"00e00",-- 224
x"00e00",-- 224
x"00f00",-- 240
x"01100",-- 272
x"01200",-- 288
x"01100",-- 272
x"00e00",-- 224
x"00b00",-- 176
x"00800",-- 128
x"00600",-- 96
x"00500",-- 80
x"00300",-- 48
x"00000",-- 0
x"ffb00",-- -80
x"ff800",-- -128
x"ff600",-- -160
x"ff500",-- -176
x"ff400",-- -192
x"ff400",-- -192
x"ff200",-- -224
x"ff000",-- -256
x"ff000",-- -256
x"ff100",-- -240
x"ff400",-- -192
x"ff600",-- -160
x"ff800",-- -128
x"ff900",-- -112
x"ffa00",-- -96
x"ffd00",-- -48
x"00000",-- 0
x"00300",-- 48
x"00600",-- 96
x"00800",-- 128
x"00900",-- 144
x"00a00",-- 160
x"00b00",-- 176
x"00d00",-- 208
x"00d00",-- 208
x"00e00",-- 224
x"00d00",-- 208
x"00c00",-- 192
x"00a00",-- 160
x"00900",-- 144
x"00900",-- 144
x"00800",-- 128
x"00600",-- 96
x"00300",-- 48
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffb00",-- -80
x"ff900",-- -112
x"ff700",-- -144
x"ff600",-- -160
x"ff600",-- -160
x"ff700",-- -144
x"ff700",-- -144
x"ff700",-- -144
x"ff700",-- -144
x"ff700",-- -144
x"ff900",-- -112
x"ffb00",-- -80
x"ffd00",-- -48
x"ffe00",-- -32
x"fff00",-- -16
x"00100",-- 16
x"00300",-- 48
x"00500",-- 80
x"00700",-- 112
x"00800",-- 128
x"00900",-- 144
x"00800",-- 128
x"00900",-- 144
x"00900",-- 144
x"00a00",-- 160
x"00900",-- 144
x"00800",-- 128
x"00700",-- 112
x"00600",-- 96
x"00400",-- 64
x"00400",-- 64
x"00300",-- 48
x"00200",-- 32
x"00000",-- 0
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffc00",-- -64
x"ffb00",-- -80
x"ffa00",-- -96
x"ff900",-- -112
x"ff900",-- -112
x"ff900",-- -112
x"ffa00",-- -96
x"ffa00",-- -96
x"ffa00",-- -96
x"ffb00",-- -80
x"ffb00",-- -80
x"ffc00",-- -64
x"ffd00",-- -48
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00300",-- 48
x"00300",-- 48
x"00500",-- 80
x"00600",-- 96
x"00600",-- 96
x"00600",-- 96
x"00600",-- 96
x"00600",-- 96
x"00500",-- 80
x"00600",-- 96
x"00500",-- 80
x"00300",-- 48
x"00200",-- 32
x"00100",-- 16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffc00",-- -64
x"ffb00",-- -80
x"ffb00",-- -80
x"ffa00",-- -96
x"ffa00",-- -96
x"ffb00",-- -80
x"ffa00",-- -96
x"ffa00",-- -96
x"ffb00",-- -80
x"ffc00",-- -64
x"ffd00",-- -48
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00300",-- 48
x"00300",-- 48
x"00400",-- 64
x"00500",-- 80
x"00500",-- 80
x"00500",-- 80
x"00500",-- 80
x"00500",-- 80
x"00500",-- 80
x"00500",-- 80
x"00400",-- 64
x"00300",-- 48
x"00300",-- 48
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffc00",-- -64
x"ffc00",-- -64
x"ffc00",-- -64
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00300",-- 48
x"00300",-- 48
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00300",-- 48
x"00300",-- 48
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00300",-- 48
x"00300",-- 48
x"00200",-- 32
x"00300",-- 48
x"00200",-- 32
x"00300",-- 48
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffc00",-- -64
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00300",-- 48
x"00300",-- 48
x"00300",-- 48
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00100",-- 16
x"fff00",-- -16
x"ffc00",-- -64
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"ffd00",-- -48
x"ffc00",-- -64
x"ffa00",-- -96
x"ffc00",-- -64
x"ffe00",-- -32
x"ffc00",-- -64
x"ff700",-- -144
x"ff400",-- -192
x"ff800",-- -128
x"ffc00",-- -64
x"ffa00",-- -96
x"ff600",-- -160
x"ff300",-- -208
x"ff200",-- -224
x"ff200",-- -224
x"fef00",-- -272
x"fef00",-- -272
x"fea00",-- -352
x"fec00",-- -320
x"fef00",-- -272
x"fee00",-- -288
x"fea00",-- -352
x"fe700",-- -400
x"fed00",-- -304
x"fef00",-- -272
x"ff300",-- -208
x"ff000",-- -256
x"fee00",-- -288
x"ff100",-- -240
x"ff800",-- -128
x"00100",-- 16
x"00200",-- 32
x"ffe00",-- -32
x"00100",-- 16
x"00500",-- 80
x"00e00",-- 224
x"01300",-- 304
x"01600",-- 352
x"01700",-- 368
x"01700",-- 368
x"02000",-- 512
x"02200",-- 544
x"02800",-- 640
x"02700",-- 624
x"02b00",-- 688
x"03000",-- 768
x"03500",-- 848
x"03b00",-- 944
x"04200",-- 1056
x"04700",-- 1136
x"05000",-- 1280
x"05000",-- 1280
x"05000",-- 1280
x"05400",-- 1344
x"05c00",-- 1472
x"05f00",-- 1520
x"05a00",-- 1440
x"05700",-- 1392
x"03800",-- 896
x"02e00",-- 736
x"03000",-- 768
x"03b00",-- 944
x"02a00",-- 672
x"00900",-- 144
x"ff200",-- -224
x"fdc00",-- -576
x"fdc00",-- -576
x"fd900",-- -624
x"fce00",-- -800
x"faf00",-- -1296
x"f9a00",-- -1632
x"f9600",-- -1696
x"f9800",-- -1664
x"f9b00",-- -1616
x"fa200",-- -1504
x"fa100",-- -1520
x"fa100",-- -1520
x"fa800",-- -1408
x"fba00",-- -1120
x"fcc00",-- -832
x"fdb00",-- -592
x"fef00",-- -272
x"ffd00",-- -48
x"00800",-- 128
x"00e00",-- 224
x"01e00",-- 480
x"02d00",-- 720
x"03700",-- 880
x"03e00",-- 992
x"03d00",-- 976
x"03500",-- 848
x"02d00",-- 720
x"03000",-- 768
x"02e00",-- 736
x"02400",-- 576
x"01500",-- 336
x"00400",-- 64
x"ff100",-- -240
x"fe500",-- -432
x"fe000",-- -512
x"fd600",-- -672
x"fc600",-- -928
x"fbb00",-- -1104
x"fad00",-- -1328
x"fa300",-- -1488
x"fa300",-- -1488
x"faa00",-- -1376
x"fad00",-- -1328
x"fa900",-- -1392
x"fa800",-- -1408
x"fad00",-- -1328
x"fba00",-- -1120
x"fd000",-- -768
x"fde00",-- -544
x"fe400",-- -448
x"fea00",-- -352
x"ff700",-- -144
x"00600",-- 96
x"01300",-- 304
x"02500",-- 592
x"02d00",-- 720
x"02f00",-- 752
x"03000",-- 768
x"03500",-- 848
x"03b00",-- 944
x"03b00",-- 944
x"03c00",-- 960
x"03400",-- 832
x"02900",-- 656
x"02000",-- 512
x"01c00",-- 448
x"01800",-- 384
x"00f00",-- 240
x"00400",-- 64
x"ff800",-- -128
x"fec00",-- -320
x"fe600",-- -416
x"fe300",-- -464
x"fde00",-- -544
x"fd700",-- -656
x"fd300",-- -720
x"fd400",-- -704
x"fd400",-- -704
x"fd600",-- -672
x"fda00",-- -608
x"fde00",-- -544
x"fe600",-- -416
x"fee00",-- -288
x"ff300",-- -208
x"ff900",-- -112
x"fff00",-- -16
x"00a00",-- 160
x"01100",-- 272
x"01700",-- 368
x"01b00",-- 432
x"01c00",-- 448
x"01e00",-- 480
x"02100",-- 528
x"02600",-- 608
x"02500",-- 592
x"01f00",-- 496
x"01a00",-- 416
x"01500",-- 336
x"01500",-- 336
x"01100",-- 272
x"00b00",-- 176
x"00300",-- 48
x"ffb00",-- -80
x"ff800",-- -128
x"ff100",-- -240
x"fef00",-- -272
x"fec00",-- -320
x"feb00",-- -336
x"fea00",-- -352
x"fe300",-- -464
x"fe700",-- -400
x"fe600",-- -416
x"fed00",-- -304
x"fee00",-- -288
x"ff200",-- -224
x"ff600",-- -160
x"ff900",-- -112
x"00400",-- 64
x"00400",-- 64
x"00b00",-- 176
x"00f00",-- 240
x"01200",-- 288
x"01600",-- 352
x"01c00",-- 448
x"02000",-- 512
x"01d00",-- 464
x"02000",-- 512
x"02300",-- 560
x"02400",-- 576
x"02600",-- 608
x"02200",-- 544
x"02200",-- 544
x"01e00",-- 480
x"01e00",-- 480
x"02100",-- 528
x"01d00",-- 464
x"02000",-- 512
x"01100",-- 272
x"01a00",-- 416
x"01e00",-- 480
x"01f00",-- 496
x"02200",-- 544
x"02300",-- 560
x"02c00",-- 704
x"02f00",-- 752
x"04100",-- 1040
x"04800",-- 1152
x"04900",-- 1168
x"04300",-- 1072
x"05400",-- 1344
x"05c00",-- 1472
x"07400",-- 1856
x"07e00",-- 2016
x"08b00",-- 2224
x"06d00",-- 1744
x"02800",-- 640
x"02600",-- 608
x"03800",-- 896
x"06900",-- 1680
x"04a00",-- 1184
x"00d00",-- 208
x"fd200",-- -736
x"fb600",-- -1184
x"fca00",-- -864
x"fd700",-- -656
x"fc700",-- -912
x"f8700",-- -1936
x"f5b00",-- -2640
x"f5b00",-- -2640
x"f7000",-- -2304
x"f7b00",-- -2128
x"f7d00",-- -2096
x"f6f00",-- -2320
x"f7100",-- -2288
x"f8200",-- -2016
x"fa100",-- -1520
x"fb600",-- -1184
x"fc300",-- -976
x"fdf00",-- -528
x"ff400",-- -192
x"00800",-- 128
x"00f00",-- 240
x"01800",-- 384
x"01d00",-- 464
x"02e00",-- 736
x"03f00",-- 1008
x"03a00",-- 928
x"02300",-- 560
x"01000",-- 256
x"00800",-- 128
x"00800",-- 128
x"00300",-- 48
x"fef00",-- -272
x"fcc00",-- -832
x"fac00",-- -1344
x"fa000",-- -1536
x"f9f00",-- -1552
x"f9800",-- -1664
x"f8900",-- -1904
x"f7a00",-- -2144
x"f6f00",-- -2320
x"f7000",-- -2304
x"f7900",-- -2160
x"f8600",-- -1952
x"f8e00",-- -1824
x"f9a00",-- -1632
x"fac00",-- -1344
x"fbe00",-- -1056
x"fce00",-- -800
x"fe200",-- -480
x"ff700",-- -144
x"01000",-- 256
x"02700",-- 624
x"03800",-- 896
x"04500",-- 1104
x"04b00",-- 1200
x"05d00",-- 1488
x"06d00",-- 1744
x"07b00",-- 1968
x"07e00",-- 2016
x"08000",-- 2048
x"08500",-- 2128
x"08b00",-- 2224
x"09600",-- 2400
x"09e00",-- 2528
x"09e00",-- 2528
x"09900",-- 2448
x"0a100",-- 2576
x"0a900",-- 2704
x"0bb00",-- 2992
x"0bc00",-- 3008
x"0c700",-- 3184
x"0a800",-- 2688
x"08e00",-- 2272
x"09400",-- 2368
x"07e00",-- 2016
x"06900",-- 1680
x"02400",-- 576
x"00300",-- 48
x"00100",-- 16
x"00400",-- 64
x"ff300",-- -208
x"fad00",-- -1328
x"f6900",-- -2416
x"f3e00",-- -3104
x"f4400",-- -3008
x"f5700",-- -2704
x"f4a00",-- -2912
x"f2300",-- -3536
x"f0600",-- -4000
x"f0e00",-- -3872
x"f3800",-- -3200
x"f5e00",-- -2592
x"f7700",-- -2192
x"f8300",-- -2000
x"f9600",-- -1696
x"fc700",-- -912
x"ffb00",-- -80
x"02300",-- 560
x"03b00",-- 944
x"05500",-- 1360
x"06f00",-- 1776
x"08b00",-- 2224
x"09400",-- 2368
x"08f00",-- 2288
x"08500",-- 2128
x"08300",-- 2096
x"08200",-- 2080
x"06d00",-- 1744
x"03e00",-- 992
x"01400",-- 320
x"00100",-- 16
x"fea00",-- -352
x"fd200",-- -736
x"fa300",-- -1488
x"f7400",-- -2240
x"f5000",-- -2816
x"f3f00",-- -3088
x"f4300",-- -3024
x"f3800",-- -3200
x"f2500",-- -3504
x"f1400",-- -3776
x"f1b00",-- -3664
x"f3500",-- -3248
x"f5500",-- -2736
x"f6e00",-- -2336
x"f7d00",-- -2096
x"f9100",-- -1776
x"fbc00",-- -1088
x"fe900",-- -368
x"01100",-- 272
x"02b00",-- 688
x"03e00",-- 992
x"05d00",-- 1488
x"07700",-- 1904
x"09000",-- 2304
x"09700",-- 2416
x"09700",-- 2416
x"09300",-- 2352
x"09800",-- 2432
x"09300",-- 2352
x"08600",-- 2144
x"07100",-- 1808
x"05900",-- 1424
x"04a00",-- 1184
x"03700",-- 880
x"02800",-- 640
x"00b00",-- 176
x"ff800",-- -128
x"fe700",-- -400
x"fe400",-- -448
x"fe200",-- -480
x"fdd00",-- -560
x"fe100",-- -496
x"fe900",-- -368
x"ff800",-- -128
x"00d00",-- 208
x"03200",-- 800
x"04300",-- 1072
x"06a00",-- 1696
x"08200",-- 2080
x"0a200",-- 2592
x"0bf00",-- 3056
x"0df00",-- 3568
x"10000",-- 4096
x"11800",-- 4480
x"12900",-- 4752
x"14e00",-- 5344
x"11f00",-- 4592
x"07c00",-- 1984
x"04500",-- 1104
x"07a00",-- 1952
x"0d500",-- 3408
x"0ae00",-- 2784
x"03300",-- 816
x"fa500",-- -1456
x"f2e00",-- -3360
x"f3500",-- -3248
x"f7900",-- -2160
x"f7900",-- -2160
x"f0200",-- -4064
x"e9c00",-- -5696
x"e8f00",-- -5904
x"eb100",-- -5360
x"edb00",-- -4688
x"f0200",-- -4064
x"efa00",-- -4192
x"ef300",-- -4304
x"f2d00",-- -3376
x"f8100",-- -2032
x"fb700",-- -1168
x"fc600",-- -928
x"ff000",-- -256
x"02800",-- 640
x"06100",-- 1552
x"08700",-- 2160
x"0a000",-- 2560
x"09000",-- 2304
x"08900",-- 2192
x"0a700",-- 2672
x"0b400",-- 2880
x"0a300",-- 2608
x"07700",-- 1904
x"04200",-- 1056
x"01900",-- 400
x"00000",-- 0
x"ff500",-- -176
x"fce00",-- -800
x"f8900",-- -1904
x"f5c00",-- -2624
x"f4100",-- -3056
x"f3100",-- -3312
x"f2200",-- -3552
x"f1700",-- -3728
x"f0800",-- -3968
x"f0300",-- -4048
x"f1c00",-- -3648
x"f3900",-- -3184
x"f4400",-- -3008
x"f5600",-- -2720
x"f7c00",-- -2112
x"faa00",-- -1376
x"fde00",-- -544
x"00600",-- 96
x"02000",-- 512
x"02d00",-- 720
x"05100",-- 1296
x"08300",-- 2096
x"0a400",-- 2624
x"0aa00",-- 2720
x"0a800",-- 2688
x"0a000",-- 2560
x"09f00",-- 2544
x"0a900",-- 2704
x"0ab00",-- 2736
x"0a000",-- 2560
x"08b00",-- 2224
x"08400",-- 2112
x"07e00",-- 2016
x"07600",-- 1888
x"07100",-- 1808
x"06e00",-- 1760
x"07800",-- 1920
x"08600",-- 2144
x"09100",-- 2320
x"09600",-- 2400
x"09c00",-- 2496
x"0ab00",-- 2736
x"0ce00",-- 3296
x"0ef00",-- 3824
x"0e600",-- 3680
x"0dc00",-- 3520
x"0b600",-- 2912
x"09800",-- 2432
x"08500",-- 2128
x"06400",-- 1600
x"05500",-- 1360
x"03300",-- 816
x"01100",-- 272
x"fe700",-- -400
x"fa800",-- -1408
x"f6500",-- -2480
x"f2300",-- -3536
x"f0e00",-- -3872
x"f0100",-- -4080
x"ef600",-- -4256
x"ede00",-- -4640
x"ec300",-- -5072
x"ebb00",-- -5200
x"ed200",-- -4832
x"efb00",-- -4176
x"f2200",-- -3552
x"f4400",-- -3008
x"f6700",-- -2448
x"f9a00",-- -1632
x"fcf00",-- -784
x"00800",-- 128
x"03c00",-- 960
x"06200",-- 1568
x"08200",-- 2080
x"09400",-- 2368
x"08900",-- 2192
x"08100",-- 2064
x"09400",-- 2368
x"0a600",-- 2656
x"09d00",-- 2512
x"06e00",-- 1760
x"03b00",-- 944
x"00900",-- 144
x"fea00",-- -352
x"fd700",-- -656
x"faf00",-- -1296
x"f7600",-- -2208
x"f4400",-- -3008
x"f2700",-- -3472
x"f1100",-- -3824
x"f0100",-- -4080
x"ef000",-- -4352
x"ee600",-- -4512
x"ee100",-- -4592
x"efa00",-- -4192
x"f1b00",-- -3664
x"f3000",-- -3328
x"f4800",-- -2944
x"f6800",-- -2432
x"f9b00",-- -1616
x"fc900",-- -880
x"ff700",-- -144
x"01e00",-- 480
x"03c00",-- 960
x"05900",-- 1424
x"08100",-- 2064
x"09d00",-- 2512
x"0b100",-- 2832
x"0bc00",-- 3008
x"0bd00",-- 3024
x"0c100",-- 3088
x"0b600",-- 2912
x"0af00",-- 2800
x"09a00",-- 2464
x"08700",-- 2160
x"07b00",-- 1968
x"07600",-- 1888
x"06900",-- 1680
x"05300",-- 1328
x"04700",-- 1136
x"03700",-- 880
x"03900",-- 912
x"04900",-- 1168
x"06300",-- 1584
x"06f00",-- 1776
x"07c00",-- 1984
x"08c00",-- 2240
x"0a500",-- 2640
x"0c800",-- 3200
x"0f200",-- 3872
x"10d00",-- 4304
x"10100",-- 4112
x"10900",-- 4240
x"0e900",-- 3728
x"0cd00",-- 3280
x"0ad00",-- 2768
x"08d00",-- 2256
x"07300",-- 1840
x"04b00",-- 1200
x"03800",-- 896
x"ffc00",-- -64
x"fae00",-- -1312
x"f5f00",-- -2576
x"f3200",-- -3296
x"f1000",-- -3840
x"efa00",-- -4192
x"ee800",-- -4480
x"ec700",-- -5008
x"eaa00",-- -5472
x"ea400",-- -5568
x"ec400",-- -5056
x"edd00",-- -4656
x"f0500",-- -4016
x"f2800",-- -3456
x"f5600",-- -2720
x"f8600",-- -1952
x"fbb00",-- -1104
x"ff700",-- -144
x"02000",-- 512
x"04700",-- 1136
x"05d00",-- 1488
x"07100",-- 1808
x"08e00",-- 2272
x"0ac00",-- 2752
x"0af00",-- 2800
x"09d00",-- 2512
x"07c00",-- 1984
x"06600",-- 1632
x"05900",-- 1424
x"03c00",-- 960
x"01500",-- 336
x"fd600",-- -672
x"fa200",-- -1504
x"f7d00",-- -2096
x"f5f00",-- -2576
x"f4200",-- -3040
x"f1900",-- -3696
x"ef800",-- -4224
x"ee700",-- -4496
x"ee900",-- -4464
x"ef400",-- -4288
x"f0000",-- -4096
x"f0b00",-- -3920
x"f2000",-- -3584
x"f4800",-- -2944
x"f7500",-- -2224
x"fa000",-- -1536
x"fc000",-- -1024
x"fe700",-- -400
x"01200",-- 288
x"03f00",-- 1008
x"06b00",-- 1712
x"08500",-- 2128
x"09700",-- 2416
x"0aa00",-- 2720
x"0bf00",-- 3056
x"0cb00",-- 3248
x"0cb00",-- 3248
x"0c200",-- 3104
x"0b400",-- 2880
x"0a700",-- 2672
x"09e00",-- 2528
x"09600",-- 2400
x"08900",-- 2192
x"07900",-- 1936
x"06f00",-- 1776
x"05e00",-- 1504
x"06200",-- 1568
x"06f00",-- 1776
x"08200",-- 2080
x"08300",-- 2096
x"08b00",-- 2224
x"0a100",-- 2576
x"0af00",-- 2800
x"0e200",-- 3616
x"0f400",-- 3904
x"0ff00",-- 4080
x"0fc00",-- 4032
x"11c00",-- 4544
x"13700",-- 4976
x"10500",-- 4176
x"0c400",-- 3136
x"08d00",-- 2256
x"06f00",-- 1776
x"05900",-- 1424
x"05300",-- 1328
x"03100",-- 784
x"fd900",-- -624
x"f7300",-- -2256
x"f3d00",-- -3120
x"f1700",-- -3728
x"ef100",-- -4336
x"ed300",-- -4816
x"eb400",-- -5312
x"e9e00",-- -5664
x"e9000",-- -5888
x"ea600",-- -5536
x"eb100",-- -5360
x"eb500",-- -5296
x"ed600",-- -4768
x"f1500",-- -3760
x"f5700",-- -2704
x"f9200",-- -1760
x"fc700",-- -912
x"fea00",-- -352
x"00700",-- 112
x"02900",-- 656
x"05b00",-- 1456
x"08800",-- 2176
x"0a700",-- 2672
x"0b200",-- 2848
x"09f00",-- 2544
x"08500",-- 2128
x"07300",-- 1840
x"06900",-- 1680
x"04c00",-- 1216
x"02800",-- 640
x"ffd00",-- -48
x"fcb00",-- -848
x"f9b00",-- -1616
x"f7000",-- -2304
x"f4900",-- -2928
x"f2100",-- -3568
x"f0500",-- -4016
x"ef800",-- -4224
x"eed00",-- -4400
x"edd00",-- -4656
x"edd00",-- -4656
x"ee600",-- -4512
x"efc00",-- -4160
x"f2300",-- -3536
x"f4c00",-- -2880
x"f6b00",-- -2384
x"f8e00",-- -1824
x"fbb00",-- -1104
x"fe800",-- -384
x"01300",-- 304
x"04000",-- 1024
x"06600",-- 1632
x"08800",-- 2176
x"0a900",-- 2704
x"0bf00",-- 3056
x"0ce00",-- 3296
x"0cd00",-- 3280
x"0d100",-- 3344
x"0d300",-- 3376
x"0ce00",-- 3296
x"0cc00",-- 3264
x"0bc00",-- 3008
x"0a800",-- 2688
x"09700",-- 2416
x"08600",-- 2144
x"07900",-- 1936
x"07900",-- 1936
x"08600",-- 2144
x"08a00",-- 2208
x"08900",-- 2192
x"08c00",-- 2240
x"08b00",-- 2224
x"09d00",-- 2512
x"0ba00",-- 2976
x"0df00",-- 3568
x"10200",-- 4128
x"10d00",-- 4304
x"10400",-- 4160
x"11e00",-- 4576
x"12500",-- 4688
x"11400",-- 4416
x"0d800",-- 3456
x"0a400",-- 2624
x"08200",-- 2080
x"05d00",-- 1488
x"05400",-- 1344
x"03a00",-- 928
x"ff300",-- -208
x"f8e00",-- -1824
x"f5800",-- -2688
x"f2500",-- -3504
x"efc00",-- -4160
x"ed800",-- -4736
x"ebb00",-- -5200
x"e9f00",-- -5648
x"e8800",-- -6016
x"ea100",-- -5616
x"ea500",-- -5552
x"eaa00",-- -5472
x"ebb00",-- -5200
x"eea00",-- -4448
x"f2100",-- -3568
x"f5a00",-- -2656
x"f9900",-- -1648
x"fbd00",-- -1072
x"fc700",-- -912
x"ff100",-- -240
x"03500",-- 848
x"05e00",-- 1504
x"08100",-- 2064
x"08600",-- 2144
x"08200",-- 2080
x"07700",-- 1904
x"07500",-- 1872
x"07300",-- 1840
x"04f00",-- 1264
x"02800",-- 640
x"01500",-- 336
x"ff600",-- -160
x"fd000",-- -768
x"fa700",-- -1424
x"f7500",-- -2224
x"f4700",-- -2960
x"f2800",-- -3456
x"f2600",-- -3488
x"f1800",-- -3712
x"f0200",-- -4064
x"ef800",-- -4224
x"efb00",-- -4176
x"f0300",-- -4048
x"f2000",-- -3584
x"f4000",-- -3072
x"f5a00",-- -2656
x"f7600",-- -2208
x"fa000",-- -1536
x"fcf00",-- -784
x"fec00",-- -320
x"01400",-- 320
x"03a00",-- 928
x"05b00",-- 1456
x"08500",-- 2128
x"0a300",-- 2608
x"0b500",-- 2896
x"0b700",-- 2928
x"0bb00",-- 2992
x"0c400",-- 3136
x"0cd00",-- 3280
x"0d500",-- 3408
x"0d500",-- 3408
x"0c800",-- 3200
x"0b600",-- 2912
x"0ac00",-- 2752
x"0a300",-- 2608
x"0a000",-- 2560
x"0a900",-- 2704
x"0ae00",-- 2784
x"0a800",-- 2688
x"0a400",-- 2624
x"0a400",-- 2624
x"0b500",-- 2896
x"0c700",-- 3184
x"0e800",-- 3712
x"10400",-- 4160
x"10900",-- 4240
x"10300",-- 4144
x"10100",-- 4112
x"11000",-- 4352
x"11000",-- 4352
x"0e500",-- 3664
x"0b700",-- 2928
x"09300",-- 2352
x"07a00",-- 1952
x"05b00",-- 1456
x"03600",-- 864
x"00500",-- 80
x"fbe00",-- -1056
x"f8c00",-- -1856
x"f6400",-- -2496
x"f3300",-- -3280
x"efb00",-- -4176
x"ece00",-- -4896
x"eb600",-- -5280
x"ea100",-- -5616
x"ea200",-- -5600
x"ea900",-- -5488
x"ea800",-- -5504
x"ea700",-- -5520
x"ec600",-- -5024
x"eef00",-- -4368
x"f1700",-- -3728
x"f3b00",-- -3152
x"f5d00",-- -2608
x"f8900",-- -1904
x"fb900",-- -1136
x"ff200",-- -224
x"01300",-- 304
x"02200",-- 544
x"03100",-- 784
x"04700",-- 1136
x"05700",-- 1392
x"06400",-- 1600
x"05f00",-- 1520
x"04600",-- 1120
x"03100",-- 784
x"02400",-- 576
x"01c00",-- 448
x"fff00",-- -16
x"fd800",-- -640
x"fb300",-- -1232
x"f9000",-- -1792
x"f7b00",-- -2128
x"f6700",-- -2448
x"f5000",-- -2816
x"f3100",-- -3312
x"f2700",-- -3472
x"f2800",-- -3456
x"f3100",-- -3312
x"f3400",-- -3264
x"f3d00",-- -3120
x"f4700",-- -2960
x"f5800",-- -2688
x"f8000",-- -2048
x"fa000",-- -1536
x"fc100",-- -1008
x"fd900",-- -624
x"ffe00",-- -32
x"02100",-- 528
x"04400",-- 1088
x"06700",-- 1648
x"07c00",-- 1984
x"09100",-- 2320
x"0a600",-- 2656
x"0bd00",-- 3024
x"0cc00",-- 3264
x"0d600",-- 3424
x"0d800",-- 3456
x"0d900",-- 3472
x"0d600",-- 3424
x"0d400",-- 3392
x"0cf00",-- 3312
x"0c800",-- 3200
x"0c300",-- 3120
x"0b800",-- 2944
x"0b500",-- 2896
x"0a600",-- 2656
x"0af00",-- 2800
x"0ae00",-- 2784
x"0b900",-- 2960
x"0c600",-- 3168
x"0c200",-- 3104
x"0d600",-- 3424
x"0d900",-- 3472
x"0dc00",-- 3520
x"0e400",-- 3648
x"0e800",-- 3712
x"0e200",-- 3616
x"0ce00",-- 3296
x"0a900",-- 2704
x"09100",-- 2320
x"07c00",-- 1984
x"06100",-- 1552
x"04d00",-- 1232
x"02200",-- 544
x"00300",-- 48
x"fd700",-- -656
x"fab00",-- -1360
x"f8400",-- -1984
x"f4800",-- -2944
x"f1b00",-- -3664
x"ef900",-- -4208
x"eeb00",-- -4432
x"ee400",-- -4544
x"ed900",-- -4720
x"ecc00",-- -4928
x"ec500",-- -5040
x"ebe00",-- -5152
x"ed400",-- -4800
x"eea00",-- -4448
x"efa00",-- -4192
x"f2500",-- -3504
x"f4500",-- -2992
x"f6f00",-- -2320
x"f8d00",-- -1840
x"fa400",-- -1472
x"fbb00",-- -1104
x"fcc00",-- -832
x"fe900",-- -368
x"00a00",-- 160
x"01600",-- 352
x"02200",-- 544
x"02500",-- 592
x"02300",-- 560
x"02600",-- 608
x"01a00",-- 416
x"01600",-- 352
x"00100",-- 16
x"ff200",-- -224
x"fe600",-- -416
x"fd100",-- -752
x"fbe00",-- -1056
x"faa00",-- -1376
x"f9800",-- -1664
x"f8e00",-- -1824
x"f8a00",-- -1888
x"f8800",-- -1920
x"f8900",-- -1904
x"f8100",-- -2032
x"f8a00",-- -1888
x"f9100",-- -1776
x"f9f00",-- -1552
x"fb600",-- -1184
x"fc700",-- -912
x"fde00",-- -544
x"ff500",-- -176
x"00d00",-- 208
x"02500",-- 592
x"03900",-- 912
x"04900",-- 1168
x"06000",-- 1536
x"06b00",-- 1712
x"07d00",-- 2000
x"08900",-- 2192
x"09000",-- 2304
x"09400",-- 2368
x"09000",-- 2304
x"09300",-- 2352
x"09200",-- 2336
x"08e00",-- 2272
x"08f00",-- 2288
x"08c00",-- 2240
x"07f00",-- 2032
x"08000",-- 2048
x"07900",-- 1936
x"07400",-- 1856
x"07a00",-- 1952
x"07e00",-- 2016
x"08400",-- 2112
x"08600",-- 2144
x"08b00",-- 2224
x"09600",-- 2400
x"0a200",-- 2592
x"0a500",-- 2640
x"0ae00",-- 2784
x"0ab00",-- 2736
x"0ae00",-- 2784
x"0b000",-- 2816
x"0a400",-- 2624
x"09d00",-- 2512
x"08e00",-- 2272
x"08a00",-- 2208
x"07800",-- 1920
x"06800",-- 1664
x"05900",-- 1424
x"04000",-- 1024
x"02300",-- 560
x"00900",-- 144
x"fef00",-- -272
x"fcd00",-- -816
x"fb300",-- -1232
x"f9700",-- -1680
x"f8500",-- -1968
x"f6900",-- -2416
x"f5800",-- -2688
x"f4900",-- -2928
x"f3500",-- -3248
x"f2c00",-- -3392
x"f2800",-- -3456
x"f2000",-- -3584
x"f1f00",-- -3600
x"f2900",-- -3440
x"f3500",-- -3248
x"f4500",-- -2992
x"f4f00",-- -2832
x"f6300",-- -2512
x"f6c00",-- -2368
x"f7c00",-- -2112
x"f9000",-- -1792
x"f9e00",-- -1568
x"fab00",-- -1360
x"fbc00",-- -1088
x"fcb00",-- -848
x"fd500",-- -688
x"fdc00",-- -576
x"fdf00",-- -528
x"fe100",-- -496
x"fd900",-- -624
x"fda00",-- -608
x"fd900",-- -624
x"fd300",-- -720
x"fd000",-- -768
x"fcd00",-- -816
x"fc800",-- -896
x"fc300",-- -976
x"fc000",-- -1024
x"fbf00",-- -1040
x"fbf00",-- -1040
x"fc200",-- -992
x"fc700",-- -912
x"fc600",-- -928
x"fc900",-- -880
x"fcd00",-- -816
x"fd200",-- -736
x"fdc00",-- -576
x"fe400",-- -448
x"ff000",-- -256
x"ff900",-- -112
x"00300",-- 48
x"00e00",-- 224
x"01300",-- 304
x"01c00",-- 448
x"02400",-- 576
x"02a00",-- 672
x"02f00",-- 752
x"03600",-- 864
x"03b00",-- 944
x"03e00",-- 992
x"04400",-- 1088
x"04700",-- 1136
x"04c00",-- 1216
x"05200",-- 1312
x"05600",-- 1376
x"05900",-- 1424
x"05c00",-- 1472
x"06200",-- 1568
x"06a00",-- 1696
x"06d00",-- 1744
x"07100",-- 1808
x"07700",-- 1904
x"07900",-- 1936
x"07f00",-- 2032
x"08100",-- 2064
x"08500",-- 2128
x"08600",-- 2144
x"08b00",-- 2224
x"08e00",-- 2272
x"08f00",-- 2288
x"09100",-- 2320
x"08e00",-- 2272
x"08b00",-- 2224
x"08400",-- 2112
x"08200",-- 2080
x"08000",-- 2048
x"07e00",-- 2016
x"07a00",-- 1952
x"07300",-- 1840
x"06a00",-- 1696
x"05e00",-- 1504
x"04f00",-- 1264
x"03f00",-- 1008
x"02d00",-- 720
x"01c00",-- 448
x"00a00",-- 160
x"ffa00",-- -96
x"fe900",-- -368
x"fd800",-- -640
x"fc500",-- -944
x"fb300",-- -1232
x"fa400",-- -1472
x"f9600",-- -1696
x"f8a00",-- -1888
x"f8000",-- -2048
x"f7a00",-- -2144
x"f7500",-- -2224
x"f7100",-- -2288
x"f6e00",-- -2336
x"f6d00",-- -2352
x"f6a00",-- -2400
x"f6d00",-- -2352
x"f6e00",-- -2336
x"f7300",-- -2256
x"f7a00",-- -2144
x"f7f00",-- -2064
x"f8600",-- -1952
x"f8800",-- -1920
x"f8800",-- -1920
x"f8600",-- -1952
x"f8700",-- -1936
x"f8700",-- -1936
x"f8700",-- -1936
x"f8a00",-- -1888
x"f8d00",-- -1840
x"f9000",-- -1792
x"f9500",-- -1712
x"f9a00",-- -1632
x"f9e00",-- -1568
x"fa300",-- -1488
x"fa800",-- -1408
x"fad00",-- -1328
x"fb400",-- -1216
x"fbc00",-- -1088
x"fc200",-- -992
x"fcb00",-- -848
x"fd200",-- -736
x"fdb00",-- -592
x"fe500",-- -432
x"fef00",-- -272
x"ffa00",-- -96
x"00400",-- 64
x"00d00",-- 208
x"01600",-- 352
x"01d00",-- 464
x"02400",-- 576
x"02a00",-- 672
x"03100",-- 784
x"03700",-- 880
x"03c00",-- 960
x"04200",-- 1056
x"04700",-- 1136
x"04c00",-- 1216
x"05000",-- 1280
x"05400",-- 1344
x"05800",-- 1408
x"05c00",-- 1472
x"05f00",-- 1520
x"06200",-- 1568
x"06600",-- 1632
x"06900",-- 1680
x"06b00",-- 1712
x"06d00",-- 1744
x"06e00",-- 1760
x"06f00",-- 1776
x"07000",-- 1792
x"07000",-- 1792
x"07000",-- 1792
x"07000",-- 1792
x"06f00",-- 1776
x"07000",-- 1792
x"07000",-- 1792
x"07000",-- 1792
x"07100",-- 1808
x"07000",-- 1792
x"06f00",-- 1776
x"06e00",-- 1760
x"06c00",-- 1728
x"06b00",-- 1712
x"06b00",-- 1712
x"06a00",-- 1696
x"06600",-- 1632
x"06100",-- 1552
x"05c00",-- 1472
x"05700",-- 1392
x"04e00",-- 1248
x"04500",-- 1104
x"03800",-- 896
x"02800",-- 640
x"01800",-- 384
x"00700",-- 112
x"ff800",-- -128
x"fe800",-- -384
x"fdb00",-- -592
x"fcf00",-- -784
x"fc400",-- -960
x"fb900",-- -1136
x"fae00",-- -1312
x"fa300",-- -1488
x"f9800",-- -1664
x"f9200",-- -1760
x"f8e00",-- -1824
x"f8c00",-- -1856
x"f8b00",-- -1872
x"f8b00",-- -1872
x"f8900",-- -1904
x"f8700",-- -1936
x"f8400",-- -1984
x"f8300",-- -2000
x"f8200",-- -2016
x"f8100",-- -2032
x"f8400",-- -1984
x"f8600",-- -1952
x"f8900",-- -1904
x"f8b00",-- -1872
x"f8b00",-- -1872
x"f8b00",-- -1872
x"f8c00",-- -1856
x"f8e00",-- -1824
x"f9000",-- -1792
x"f9400",-- -1728
x"f9900",-- -1648
x"f9e00",-- -1568
x"fa400",-- -1472
x"fac00",-- -1344
x"fb200",-- -1248
x"fb700",-- -1168
x"fbe00",-- -1056
x"fc700",-- -912
x"fcf00",-- -784
x"fd800",-- -640
x"fe100",-- -496
x"fe900",-- -368
x"ff100",-- -240
x"ffa00",-- -96
x"00200",-- 32
x"00900",-- 144
x"00f00",-- 240
x"01500",-- 336
x"01b00",-- 432
x"02100",-- 528
x"02700",-- 624
x"02c00",-- 704
x"03100",-- 784
x"03600",-- 864
x"03b00",-- 944
x"03f00",-- 1008
x"04300",-- 1072
x"04500",-- 1104
x"04600",-- 1120
x"04600",-- 1120
x"04600",-- 1120
x"04800",-- 1152
x"04800",-- 1152
x"04700",-- 1136
x"04700",-- 1136
x"04700",-- 1136
x"04700",-- 1136
x"04700",-- 1136
x"04600",-- 1120
x"04500",-- 1104
x"04400",-- 1088
x"04400",-- 1088
x"04500",-- 1104
x"04500",-- 1104
x"04600",-- 1120
x"04600",-- 1120
x"04600",-- 1120
x"04500",-- 1104
x"04500",-- 1104
x"04400",-- 1088
x"04200",-- 1056
x"04100",-- 1040
x"04000",-- 1024
x"03e00",-- 992
x"03b00",-- 944
x"03800",-- 896
x"03500",-- 848
x"03300",-- 816
x"03000",-- 768
x"02e00",-- 736
x"02c00",-- 704
x"02a00",-- 672
x"02800",-- 640
x"02500",-- 592
x"02300",-- 560
x"01f00",-- 496
x"01c00",-- 448
x"01700",-- 368
x"01200",-- 288
x"00c00",-- 192
x"00700",-- 112
x"00100",-- 16
x"ffb00",-- -80
x"ff500",-- -176
x"fef00",-- -272
x"fea00",-- -352
x"fe500",-- -432
x"fe000",-- -512
x"fdc00",-- -576
x"fd900",-- -624
x"fd600",-- -672
x"fd300",-- -720
x"fd100",-- -752
x"fce00",-- -800
x"fcc00",-- -832
x"fc900",-- -880
x"fc600",-- -928
x"fc300",-- -976
x"fc100",-- -1008
x"fbf00",-- -1040
x"fbc00",-- -1088
x"fb900",-- -1136
x"fb700",-- -1168
x"fb600",-- -1184
x"fb400",-- -1216
x"fb300",-- -1232
x"fb200",-- -1248
x"fb000",-- -1280
x"fb000",-- -1280
x"fb100",-- -1264
x"fb100",-- -1264
x"fb300",-- -1232
x"fb500",-- -1200
x"fb700",-- -1168
x"fb900",-- -1136
x"fbc00",-- -1088
x"fbf00",-- -1040
x"fc300",-- -976
x"fc700",-- -912
x"fcb00",-- -848
x"fcf00",-- -784
x"fd300",-- -720
x"fd800",-- -640
x"fdc00",-- -576
x"fe200",-- -480
x"fe700",-- -400
x"feb00",-- -336
x"ff000",-- -256
x"ff500",-- -176
x"ff900",-- -112
x"ffe00",-- -32
x"00200",-- 32
x"00600",-- 96
x"00b00",-- 176
x"00f00",-- 240
x"01300",-- 304
x"01600",-- 352
x"01a00",-- 416
x"01d00",-- 464
x"02100",-- 528
x"02400",-- 576
x"02700",-- 624
x"02a00",-- 672
x"02d00",-- 720
x"02f00",-- 752
x"03100",-- 784
x"03300",-- 816
x"03500",-- 848
x"03600",-- 864
x"03700",-- 880
x"03700",-- 880
x"03700",-- 880
x"03700",-- 880
x"03700",-- 880
x"03700",-- 880
x"03600",-- 864
x"03500",-- 848
x"03400",-- 832
x"03200",-- 800
x"03100",-- 784
x"02f00",-- 752
x"02d00",-- 720
x"02a00",-- 672
x"02800",-- 640
x"02600",-- 608
x"02300",-- 560
x"02100",-- 528
x"01e00",-- 480
x"01b00",-- 432
x"01900",-- 400
x"01700",-- 368
x"01400",-- 320
x"01200",-- 288
x"01000",-- 256
x"00e00",-- 224
x"00c00",-- 192
x"00a00",-- 160
x"00900",-- 144
x"00700",-- 112
x"00500",-- 80
x"00400",-- 64
x"00300",-- 48
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"ffd00",-- -48
x"ffc00",-- -64
x"ffb00",-- -80
x"ffa00",-- -96
x"ff900",-- -112
x"ff800",-- -128
x"ff700",-- -144
x"ff500",-- -176
x"ff400",-- -192
x"ff300",-- -208
x"ff100",-- -240
x"ff000",-- -256
x"fef00",-- -272
x"fed00",-- -304
x"fec00",-- -320
x"feb00",-- -336
x"fe900",-- -368
x"fe800",-- -384
x"fe700",-- -400
x"fe600",-- -416
x"fe600",-- -416
x"fe400",-- -448
x"fe400",-- -448
x"fe300",-- -464
x"fe300",-- -464
x"fe300",-- -464
x"fe300",-- -464
x"fe300",-- -464
x"fe200",-- -480
x"fe200",-- -480
x"fe300",-- -464
x"fe200",-- -480
x"fe200",-- -480
x"fe200",-- -480
x"fe300",-- -464
x"fe300",-- -464
x"fe300",-- -464
x"fe500",-- -432
x"fe500",-- -432
x"fe500",-- -432
x"fe700",-- -400
x"fe800",-- -384
x"fe900",-- -368
x"fea00",-- -352
x"fec00",-- -320
x"fed00",-- -304
x"fef00",-- -272
x"ff100",-- -240
x"ff300",-- -208
x"ff500",-- -176
x"ff600",-- -160
x"ff800",-- -128
x"ffa00",-- -96
x"ffc00",-- -64
x"fff00",-- -16
x"00200",-- 32
x"00400",-- 64
x"00600",-- 96
x"00900",-- 144
x"00b00",-- 176
x"00e00",-- 224
x"00f00",-- 240
x"01100",-- 272
x"01300",-- 304
x"01500",-- 336
x"01600",-- 352
x"01800",-- 384
x"01900",-- 400
x"01a00",-- 416
x"01b00",-- 432
x"01b00",-- 432
x"01b00",-- 432
x"01b00",-- 432
x"01c00",-- 448
x"01c00",-- 448
x"01c00",-- 448
x"01c00",-- 448
x"01b00",-- 432
x"01b00",-- 432
x"01a00",-- 416
x"01900",-- 400
x"01900",-- 400
x"01800",-- 384
x"01600",-- 352
x"01600",-- 352
x"01500",-- 336
x"01300",-- 304
x"01300",-- 304
x"01100",-- 272
x"00f00",-- 240
x"00d00",-- 208
x"00c00",-- 192
x"00a00",-- 160
x"00900",-- 144
x"00700",-- 112
x"00500",-- 80
x"00300",-- 48
x"00100",-- 16
x"00000",-- 0
x"ffd00",-- -48
x"ffc00",-- -64
x"ffa00",-- -96
x"ff900",-- -112
x"ff700",-- -144
x"ff600",-- -160
x"ff400",-- -192
x"ff300",-- -208
x"ff200",-- -224
x"ff200",-- -224
x"ff100",-- -240
x"ff100",-- -240
x"ff000",-- -256
x"ff000",-- -256
x"fef00",-- -272
x"fef00",-- -272
x"ff000",-- -256
x"ff000",-- -256
x"ff000",-- -256
x"ff000",-- -256
x"ff000",-- -256
x"ff000",-- -256
x"ff100",-- -240
x"ff100",-- -240
x"ff200",-- -224
x"ff300",-- -208
x"ff300",-- -208
x"ff300",-- -208
x"ff400",-- -192
x"ff500",-- -176
x"ff600",-- -160
x"ff600",-- -160
x"ff700",-- -144
x"ff700",-- -144
x"ff800",-- -128
x"ff800",-- -128
x"ff900",-- -112
x"ffa00",-- -96
x"ffb00",-- -80
x"ffc00",-- -64
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00300",-- 48
x"00400",-- 64
x"00400",-- 64
x"00500",-- 80
x"00600",-- 96
x"00600",-- 96
x"00600",-- 96
x"00700",-- 112
x"00700",-- 112
x"00800",-- 128
x"00700",-- 112
x"00800",-- 128
x"00800",-- 128
x"00800",-- 128
x"00800",-- 128
x"00900",-- 144
x"00900",-- 144
x"00900",-- 144
x"00900",-- 144
x"00900",-- 144
x"00a00",-- 160
x"00a00",-- 160
x"00a00",-- 160
x"00a00",-- 160
x"00a00",-- 160
x"00a00",-- 160
x"00a00",-- 160
x"00a00",-- 160
x"00a00",-- 160
x"00900",-- 144
x"00900",-- 144
x"00900",-- 144
x"00900",-- 144
x"00800",-- 128
x"00800",-- 128
x"00700",-- 112
x"00700",-- 112
x"00700",-- 112
x"00600",-- 96
x"00600",-- 96
x"00500",-- 80
x"00400",-- 64
x"00300",-- 48
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffc00",-- -64
x"ffc00",-- -64
x"ffb00",-- -80
x"ffb00",-- -80
x"ffc00",-- -64
x"ffb00",-- -80
x"ffa00",-- -96
x"ffa00",-- -96
x"ffa00",-- -96
x"ff900",-- -112
x"ff900",-- -112
x"ff900",-- -112
x"ff800",-- -128
x"ff800",-- -128
x"ff700",-- -144
x"ff700",-- -144
x"ff600",-- -160
x"ff600",-- -160
x"ff500",-- -176
x"ff500",-- -176
x"ff500",-- -176
x"ff500",-- -176
x"ff500",-- -176
x"ff400",-- -192
x"ff400",-- -192
x"ff400",-- -192
x"ff400",-- -192
x"ff400",-- -192
x"ff500",-- -176
x"ff500",-- -176
x"ff600",-- -160
x"ff600",-- -160
x"ff700",-- -144
x"ff700",-- -144
x"ff700",-- -144
x"ff800",-- -128
x"ff900",-- -112
x"ff900",-- -112
x"ff900",-- -112
x"ffa00",-- -96
x"ffa00",-- -96
x"ffb00",-- -80
x"ffc00",-- -64
x"ffc00",-- -64
x"ffc00",-- -64
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00300",-- 48
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00500",-- 80
x"00600",-- 96
x"00700",-- 112
x"00700",-- 112
x"00700",-- 112
x"00700",-- 112
x"00700",-- 112
x"00800",-- 128
x"00900",-- 144
x"00900",-- 144
x"00900",-- 144
x"00900",-- 144
x"00900",-- 144
x"00900",-- 144
x"00900",-- 144
x"00a00",-- 160
x"00900",-- 144
x"00900",-- 144
x"00900",-- 144
x"00900",-- 144
x"00800",-- 128
x"00800",-- 128
x"00700",-- 112
x"00700",-- 112
x"00700",-- 112
x"00600",-- 96
x"00600",-- 96
x"00500",-- 80
x"00500",-- 80
x"00500",-- 80
x"00400",-- 64
x"00300",-- 48
x"00300",-- 48
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffc00",-- -64
x"ffc00",-- -64
x"ffb00",-- -80
x"ffc00",-- -64
x"ffb00",-- -80
x"ffb00",-- -80
x"ffb00",-- -80
x"ffa00",-- -96
x"ffa00",-- -96
x"ffa00",-- -96
x"ff900",-- -112
x"ff900",-- -112
x"ff900",-- -112
x"ff900",-- -112
x"ff900",-- -112
x"ff900",-- -112
x"ff900",-- -112
x"ffa00",-- -96
x"ffa00",-- -96
x"ffa00",-- -96
x"ffa00",-- -96
x"ffa00",-- -96
x"ffb00",-- -80
x"ffb00",-- -80
x"ffb00",-- -80
x"ffc00",-- -64
x"ffb00",-- -80
x"ffc00",-- -64
x"ffc00",-- -64
x"ffc00",-- -64
x"ffc00",-- -64
x"ffc00",-- -64
x"ffc00",-- -64
x"ffd00",-- -48
x"ffd00",-- -48
x"ffc00",-- -64
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00300",-- 48
x"00200",-- 32
x"00200",-- 32
x"00400",-- 64
x"00200",-- 32
x"00300",-- 48
x"00200",-- 32
x"00200",-- 32
x"00500",-- 80
x"00100",-- 16
x"00300",-- 48
x"00300",-- 48
x"00200",-- 32
x"00300",-- 48
x"00200",-- 32
x"00100",-- 16
x"00300",-- 48
x"00200",-- 32
x"00200",-- 32
x"00300",-- 48
x"00100",-- 16
x"00300",-- 48
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffd00",-- -48
x"ffe00",-- -32
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"ffd00",-- -48
x"00100",-- 16
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"ffe00",-- -32
x"00100",-- 16
x"fff00",-- -16
x"00100",-- 16
x"ffd00",-- -48
x"00100",-- 16
x"00000",-- 0
x"ffe00",-- -32
x"00100",-- 16
x"fff00",-- -16
x"00100",-- 16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00100",-- 16
x"00200",-- 32
x"fff00",-- -16
x"00200",-- 32
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"fff00",-- -16
x"00200",-- 32
x"00000",-- 0
x"00300",-- 48
x"ffe00",-- -32
x"00300",-- 48
x"00000",-- 0
x"00200",-- 32
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"00300",-- 48
x"ffe00",-- -32
x"00200",-- 32
x"00000",-- 0
x"00100",-- 16
x"fff00",-- -16
x"00200",-- 32
x"00000",-- 0
x"00400",-- 64
x"fff00",-- -16
x"ffd00",-- -48
x"00200",-- 32
x"ffa00",-- -96
x"fff00",-- -16
x"ffd00",-- -48
x"fff00",-- -16
x"ffc00",-- -64
x"ffc00",-- -64
x"ffd00",-- -48
x"ffc00",-- -64
x"ffa00",-- -96
x"ff800",-- -128
x"ffc00",-- -64
x"ffa00",-- -96
x"00300",-- 48
x"fff00",-- -16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"00500",-- 80
x"ffd00",-- -48
x"00200",-- 32
x"00300",-- 48
x"fff00",-- -16
x"00200",-- 32
x"00300",-- 48
x"00100",-- 16
x"00500",-- 80
x"fff00",-- -16
x"00000",-- 0
x"00300",-- 48
x"ffe00",-- -32
x"00300",-- 48
x"ff800",-- -128
x"ffd00",-- -48
x"00200",-- 32
x"ffa00",-- -96
x"00100",-- 16
x"00000",-- 0
x"ffb00",-- -80
x"00000",-- 0
x"fff00",-- -16
x"ff900",-- -112
x"fff00",-- -16
x"00200",-- 32
x"00200",-- 32
x"ff500",-- -176
x"00400",-- 64
x"ffc00",-- -64
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"00100",-- 16
x"ff900",-- -112
x"00600",-- 96
x"ffa00",-- -96
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"ffc00",-- -64
x"00500",-- 80
x"00500",-- 80
x"fff00",-- -16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00300",-- 48
x"ffc00",-- -64
x"00900",-- 144
x"00300",-- 48
x"fff00",-- -16
x"00300",-- 48
x"00300",-- 48
x"00000",-- 0
x"fff00",-- -16
x"00600",-- 96
x"00100",-- 16
x"00600",-- 96
x"ffa00",-- -96
x"00100",-- 16
x"00100",-- 16
x"00500",-- 80
x"00100",-- 16
x"ffa00",-- -96
x"00900",-- 144
x"ffd00",-- -48
x"00800",-- 128
x"ffd00",-- -48
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"ffd00",-- -48
x"00600",-- 96
x"00100",-- 16
x"fff00",-- -16
x"00100",-- 16
x"00000",-- 0
x"00500",-- 80
x"ffe00",-- -32
x"00900",-- 144
x"ff800",-- -128
x"00500",-- 80
x"ffd00",-- -48
x"00800",-- 128
x"ffa00",-- -96
x"00100",-- 16
x"00000",-- 0
x"ffc00",-- -64
x"00d00",-- 208
x"ff100",-- -240
x"00b00",-- 176
x"ffe00",-- -32
x"00400",-- 64
x"ffc00",-- -64
x"00100",-- 16
x"ffd00",-- -48
x"ffe00",-- -32
x"00300",-- 48
x"ff800",-- -128
x"00600",-- 96
x"ff600",-- -160
x"00500",-- 80
x"ffa00",-- -96
x"00300",-- 48
x"ff900",-- -112
x"ffe00",-- -32
x"ffd00",-- -48
x"00200",-- 32
x"00000",-- 0
x"ff400",-- -192
x"00400",-- 64
x"ffe00",-- -32
x"fff00",-- -16
x"00200",-- 32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00300",-- 48
x"ff900",-- -112
x"fff00",-- -16
x"ffb00",-- -80
x"00300",-- 48
x"ffb00",-- -80
x"00200",-- 32
x"00000",-- 0
x"ffc00",-- -64
x"00200",-- 32
x"fff00",-- -16
x"00600",-- 96
x"ffc00",-- -64
x"ffa00",-- -96
x"00500",-- 80
x"ff800",-- -128
x"00700",-- 112
x"ffc00",-- -64
x"00300",-- 48
x"ffa00",-- -96
x"fff00",-- -16
x"00300",-- 48
x"ff800",-- -128
x"00500",-- 80
x"ffe00",-- -32
x"ff900",-- -112
x"00a00",-- 160
x"ff100",-- -240
x"00900",-- 144
x"00400",-- 64
x"ff600",-- -160
x"00d00",-- 208
x"ffa00",-- -96
x"00100",-- 16
x"ffa00",-- -96
x"00000",-- 0
x"00100",-- 16
x"ffc00",-- -64
x"00300",-- 48
x"00100",-- 16
x"00400",-- 64
x"ffe00",-- -32
x"00100",-- 16
x"ffc00",-- -64
x"00000",-- 0
x"ffc00",-- -64
x"ffe00",-- -32
x"00300",-- 48
x"ffb00",-- -80
x"00100",-- 16
x"00300",-- 48
x"00400",-- 64
x"00300",-- 48
x"00200",-- 32
x"ffd00",-- -48
x"ffe00",-- -32
x"ffa00",-- -96
x"00900",-- 144
x"ffb00",-- -80
x"00800",-- 128
x"ffa00",-- -96
x"00100",-- 16
x"00400",-- 64
x"ffa00",-- -96
x"00a00",-- 160
x"ff200",-- -224
x"00f00",-- 240
x"ff500",-- -176
x"00100",-- 16
x"00700",-- 112
x"ff300",-- -208
x"00600",-- 96
x"ffe00",-- -32
x"00100",-- 16
x"ffa00",-- -96
x"00d00",-- 208
x"ff900",-- -112
x"00800",-- 128
x"ff500",-- -176
x"00500",-- 80
x"ffb00",-- -80
x"ff600",-- -160
x"00a00",-- 160
x"ff100",-- -240
x"00800",-- 128
x"ff900",-- -112
x"00a00",-- 160
x"ff600",-- -160
x"00700",-- 112
x"ff900",-- -112
x"00500",-- 80
x"fff00",-- -16
x"ff400",-- -192
x"00a00",-- 160
x"ff700",-- -144
x"00600",-- 96
x"ff800",-- -128
x"ffe00",-- -32
x"ffd00",-- -48
x"00700",-- 112
x"ff900",-- -112
x"00600",-- 96
x"fff00",-- -16
x"ff300",-- -208
x"00300",-- 48
x"00600",-- 96
x"00600",-- 96
x"ff900",-- -112
x"00900",-- 144
x"ff800",-- -128
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"00100",-- 16
x"00700",-- 112
x"ffc00",-- -64
x"fff00",-- -16
x"00600",-- 96
x"ff900",-- -112
x"00600",-- 96
x"ffc00",-- -64
x"00c00",-- 192
x"00300",-- 48
x"ff700",-- -144
x"01000",-- 256
x"fef00",-- -272
x"01100",-- 272
x"ffc00",-- -64
x"ffd00",-- -48
x"00a00",-- 160
x"ff300",-- -208
x"00800",-- 128
x"ff900",-- -112
x"00900",-- 144
x"ffe00",-- -32
x"00400",-- 64
x"00200",-- 32
x"00100",-- 16
x"ffe00",-- -32
x"ffa00",-- -96
x"00f00",-- 240
x"ffa00",-- -96
x"00400",-- 64
x"ffa00",-- -96
x"00400",-- 64
x"00200",-- 32
x"ffc00",-- -64
x"00000",-- 0
x"00600",-- 96
x"ffa00",-- -96
x"ffd00",-- -48
x"00900",-- 144
x"ffe00",-- -32
x"00900",-- 144
x"00200",-- 32
x"ffb00",-- -80
x"00600",-- 96
x"ffd00",-- -48
x"00800",-- 128
x"ffd00",-- -48
x"ffa00",-- -96
x"00600",-- 96
x"ff400",-- -192
x"00700",-- 112
x"00400",-- 64
x"fff00",-- -16
x"00a00",-- 160
x"ff900",-- -112
x"ffe00",-- -32
x"00200",-- 32
x"fff00",-- -16
x"ff900",-- -112
x"00c00",-- 192
x"ff400",-- -192
x"00b00",-- 176
x"ffc00",-- -64
x"00200",-- 32
x"00100",-- 16
x"ff400",-- -192
x"01100",-- 272
x"ff400",-- -192
x"ffe00",-- -32
x"00300",-- 48
x"ff800",-- -128
x"00500",-- 80
x"00600",-- 96
x"ff900",-- -112
x"00500",-- 80
x"ff900",-- -112
x"ffe00",-- -32
x"fff00",-- -16
x"00200",-- 32
x"00000",-- 0
x"ff800",-- -128
x"00200",-- 32
x"fff00",-- -16
x"00800",-- 128
x"ffd00",-- -48
x"fff00",-- -16
x"00600",-- 96
x"fec00",-- -320
x"00b00",-- 176
x"ffc00",-- -64
x"ff800",-- -128
x"00900",-- 144
x"ff400",-- -192
x"00100",-- 16
x"ffd00",-- -48
x"00500",-- 80
x"00d00",-- 208
x"fe800",-- -384
x"01200",-- 288
x"ff800",-- -128
x"ff200",-- -224
x"01400",-- 320
x"fee00",-- -288
x"00a00",-- 160
x"00300",-- 48
x"ffb00",-- -80
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00d00",-- 208
x"ffa00",-- -96
x"ffa00",-- -96
x"00200",-- 32
x"00000",-- 0
x"ffc00",-- -64
x"ff700",-- -144
x"00200",-- 32
x"ff700",-- -144
x"00d00",-- 208
x"ff800",-- -128
x"00e00",-- 224
x"ff200",-- -224
x"00600",-- 96
x"00400",-- 64
x"ff200",-- -224
x"01300",-- 304
x"fe900",-- -368
x"01100",-- 272
x"ff300",-- -208
x"ffe00",-- -32
x"00a00",-- 160
x"ff700",-- -144
x"00800",-- 128
x"ffc00",-- -64
x"00200",-- 32
x"00900",-- 144
x"00000",-- 0
x"ff800",-- -128
x"00b00",-- 176
x"ff600",-- -160
x"00100",-- 16
x"00700",-- 112
x"ff300",-- -208
x"01500",-- 336
x"fee00",-- -288
x"01300",-- 304
x"ff200",-- -224
x"00400",-- 64
x"00b00",-- 176
x"ff300",-- -208
x"00800",-- 128
x"ff500",-- -176
x"00000",-- 0
x"ffb00",-- -80
x"00300",-- 48
x"ffe00",-- -32
x"ffe00",-- -32
x"00800",-- 128
x"ffa00",-- -96
x"00a00",-- 160
x"ff500",-- -176
x"ff900",-- -112
x"01000",-- 256
x"fe900",-- -368
x"00b00",-- 176
x"00300",-- 48
x"feb00",-- -336
x"01900",-- 400
x"ffa00",-- -96
x"00500",-- 80
x"00c00",-- 192
x"fed00",-- -304
x"01000",-- 256
x"ff700",-- -144
x"ff700",-- -144
x"01100",-- 272
x"fee00",-- -288
x"00700",-- 112
x"00200",-- 32
x"ffc00",-- -64
x"00300",-- 48
x"ff500",-- -176
x"00500",-- 80
x"00400",-- 64
x"fff00",-- -16
x"00100",-- 16
x"00000",-- 0
x"ffd00",-- -48
x"fff00",-- -16
x"ff000",-- -256
x"ffc00",-- -64
x"01600",-- 352
x"ff500",-- -176
x"00400",-- 64
x"00000",-- 0
x"ff900",-- -112
x"00600",-- 96
x"ffe00",-- -32
x"ffc00",-- -64
x"00600",-- 96
x"fe500",-- -432
x"01300",-- 304
x"00900",-- 144
x"feb00",-- -336
x"01500",-- 336
x"ff300",-- -208
x"00a00",-- 160
x"ff400",-- -192
x"fff00",-- -16
x"00500",-- 80
x"ff900",-- -112
x"ffd00",-- -48
x"00800",-- 128
x"00300",-- 48
x"ff800",-- -128
x"00000",-- 0
x"00500",-- 80
x"ff600",-- -160
x"00400",-- 64
x"00300",-- 48
x"00100",-- 16
x"ffe00",-- -32
x"ffe00",-- -32
x"01400",-- 320
x"fe600",-- -416
x"01500",-- 336
x"feb00",-- -336
x"01000",-- 256
x"ff300",-- -208
x"ffc00",-- -64
x"01000",-- 256
x"fee00",-- -288
x"01600",-- 352
x"fe500",-- -432
x"01c00",-- 448
x"fec00",-- -320
x"00200",-- 32
x"00500",-- 80
x"fea00",-- -352
x"01800",-- 384
x"fed00",-- -304
x"00c00",-- 192
x"fee00",-- -288
x"00800",-- 128
x"ffa00",-- -96
x"00d00",-- 208
x"fed00",-- -304
x"00b00",-- 176
x"ff600",-- -160
x"ff600",-- -160
x"00700",-- 112
x"fef00",-- -272
x"02300",-- 560
x"fd800",-- -640
x"02200",-- 544
x"fe300",-- -464
x"01f00",-- 496
x"fdf00",-- -528
x"00c00",-- 192
x"00400",-- 64
x"fee00",-- -288
x"03000",-- 768
x"fc200",-- -992
x"04100",-- 1040
x"fc600",-- -928
x"01200",-- 288
x"01000",-- 256
x"fee00",-- -288
x"01400",-- 320
x"fd200",-- -736
x"02600",-- 608
x"fee00",-- -288
x"00c00",-- 192
x"ff200",-- -224
x"00f00",-- 240
x"fed00",-- -304
x"ffd00",-- -48
x"01000",-- 256
x"fe400",-- -448
x"00900",-- 144
x"ff700",-- -144
x"00d00",-- 208
x"ff800",-- -128
x"00700",-- 112
x"ff500",-- -176
x"ff800",-- -128
x"01400",-- 320
x"ff000",-- -256
x"01800",-- 384
x"fe400",-- -448
x"00c00",-- 192
x"00500",-- 80
x"ffc00",-- -64
x"00e00",-- 224
x"ff500",-- -176
x"00600",-- 96
x"fe500",-- -432
x"01b00",-- 432
x"ff100",-- -240
x"00100",-- 16
x"00900",-- 144
x"ff200",-- -224
x"01700",-- 368
x"fe400",-- -448
x"01600",-- 352
x"fef00",-- -272
x"00700",-- 112
x"00100",-- 16
x"fec00",-- -320
x"01400",-- 320
x"fef00",-- -272
x"00400",-- 64
x"01100",-- 272
x"00400",-- 64
x"fff00",-- -16
x"00300",-- 48
x"fe500",-- -432
x"01200",-- 288
x"fe900",-- -368
x"02000",-- 512
x"fe400",-- -448
x"00f00",-- 240
x"ffb00",-- -80
x"ff900",-- -112
x"01f00",-- 496
x"fea00",-- -352
x"01100",-- 272
x"fed00",-- -304
x"ff900",-- -112
x"00100",-- 16
x"00900",-- 144
x"01400",-- 320
x"ff400",-- -192
x"00d00",-- 208
x"fe200",-- -480
x"01300",-- 304
x"00100",-- 16
x"fef00",-- -272
x"01f00",-- 496
x"fd500",-- -688
x"01500",-- 336
x"fe800",-- -384
x"01c00",-- 448
x"fdc00",-- -576
x"00800",-- 128
x"01200",-- 288
x"fdd00",-- -560
x"02900",-- 656
x"fdd00",-- -560
x"02100",-- 528
x"feb00",-- -336
x"00b00",-- 176
x"00800",-- 128
x"ff200",-- -224
x"ffe00",-- -32
x"00d00",-- 208
x"00900",-- 144
x"ffa00",-- -96
x"01a00",-- 416
x"ff300",-- -208
x"ffe00",-- -32
x"00a00",-- 160
x"ffa00",-- -96
x"ffe00",-- -32
x"00a00",-- 160
x"fe700",-- -400
x"00e00",-- 224
x"fea00",-- -352
x"00700",-- 112
x"fec00",-- -320
x"fe000",-- -512
x"02b00",-- 688
x"fe000",-- -512
x"00e00",-- 224
x"00b00",-- 176
x"fed00",-- -304
x"01c00",-- 448
x"ff300",-- -208
x"fff00",-- -16
x"ffc00",-- -64
x"ff300",-- -208
x"01d00",-- 464
x"ff500",-- -176
x"ff600",-- -160
x"01c00",-- 448
x"00500",-- 80
x"00500",-- 80
x"ff900",-- -112
x"00b00",-- 176
x"ffe00",-- -32
x"ff200",-- -224
x"ffe00",-- -32
x"ff500",-- -176
x"00100",-- 16
x"00200",-- 32
x"ffd00",-- -48
x"00600",-- 96
x"00100",-- 16
x"00300",-- 48
x"00600",-- 96
x"fee00",-- -288
x"01300",-- 304
x"ff300",-- -208
x"fe100",-- -496
x"00300",-- 48
x"00400",-- 64
x"fd700",-- -656
x"01600",-- 352
x"00700",-- 112
x"fff00",-- -16
x"fea00",-- -352
x"00b00",-- 176
x"01100",-- 272
x"fde00",-- -544
x"01300",-- 304
x"ff500",-- -176
x"00000",-- 0
x"00300",-- 48
x"01300",-- 304
x"fec00",-- -320
x"01500",-- 336
x"fff00",-- -16
x"ffb00",-- -80
x"00d00",-- 208
x"00000",-- 0
x"00b00",-- 176
x"fe900",-- -368
x"00300",-- 48
x"00800",-- 128
x"ffd00",-- -48
x"ff700",-- -144
x"01e00",-- 480
x"fe400",-- -448
x"00f00",-- 240
x"ff600",-- -160
x"ff800",-- -128
x"01000",-- 256
x"fe500",-- -432
x"01b00",-- 432
x"fd500",-- -688
x"01400",-- 320
x"fed00",-- -304
x"00100",-- 16
x"ffe00",-- -32
x"ff300",-- -208
x"00d00",-- 208
x"ff100",-- -240
x"01e00",-- 480
x"fe700",-- -400
x"00500",-- 80
x"ff300",-- -208
x"02400",-- 576
x"fe200",-- -480
x"01f00",-- 496
x"00d00",-- 208
x"fed00",-- -304
x"01a00",-- 416
x"fd900",-- -624
x"01c00",-- 448
x"fe200",-- -480
x"02900",-- 656
x"ff000",-- -256
x"00d00",-- 208
x"01000",-- 256
x"fcb00",-- -848
x"03500",-- 848
x"fcc00",-- -832
x"02300",-- 560
x"00c00",-- 192
x"fe500",-- -432
x"01600",-- 352
x"fdf00",-- -528
x"00100",-- 16
x"ff700",-- -144
x"00e00",-- 224
x"ffe00",-- -32
x"ff100",-- -240
x"01400",-- 320
x"fee00",-- -288
x"00f00",-- 240
x"fe200",-- -480
x"00a00",-- 160
x"00200",-- 32
x"ff600",-- -160
x"02700",-- 624
x"ffb00",-- -80
x"ff100",-- -240
x"00900",-- 144
x"ff800",-- -128
x"01500",-- 336
x"ffa00",-- -96
x"fe800",-- -384
x"03200",-- 800
x"fd900",-- -624
x"03000",-- 768
x"fec00",-- -320
x"00300",-- 48
x"00000",-- 0
x"fdb00",-- -592
x"01500",-- 336
x"ff000",-- -256
x"00c00",-- 192
x"ff200",-- -224
x"02700",-- 624
x"fe500",-- -432
x"ff100",-- -240
x"00800",-- 128
x"ffc00",-- -64
x"00c00",-- 192
x"ff500",-- -176
x"02b00",-- 688
x"fdf00",-- -528
x"01b00",-- 432
x"ff100",-- -240
x"00000",-- 0
x"00800",-- 128
x"fda00",-- -608
x"02200",-- 544
x"fed00",-- -304
x"ffd00",-- -48
x"00e00",-- 224
x"fe800",-- -384
x"ff800",-- -128
x"00600",-- 96
x"01c00",-- 448
x"ff900",-- -112
x"ff900",-- -112
x"01f00",-- 496
x"fdc00",-- -576
x"01e00",-- 480
x"fe500",-- -432
x"00d00",-- 208
x"ff600",-- -160
x"00300",-- 48
x"01400",-- 320
x"fdb00",-- -592
x"03e00",-- 992
x"fb200",-- -1248
x"02e00",-- 736
x"ff300",-- -208
x"00100",-- 16
x"01f00",-- 496
x"00b00",-- 176
x"ff600",-- -160
x"fff00",-- -16
x"01400",-- 320
x"fc400",-- -960
x"02200",-- 544
x"fdb00",-- -592
x"03000",-- 768
x"ff800",-- -128
x"00200",-- 32
x"01000",-- 256
x"fdc00",-- -576
x"03400",-- 832
x"fcf00",-- -784
x"ffe00",-- -32
x"ffb00",-- -80
x"00a00",-- 160
x"fe900",-- -368
x"02100",-- 528
x"fed00",-- -304
x"fe400",-- -448
x"02a00",-- 672
x"fcc00",-- -832
x"04100",-- 1040
x"fc300",-- -976
x"03600",-- 864
x"fd900",-- -624
x"00900",-- 144
x"00100",-- 16
x"fda00",-- -608
x"03100",-- 784
x"fe200",-- -480
x"00100",-- 16
x"00c00",-- 192
x"01d00",-- 464
x"fc000",-- -1024
x"03d00",-- 976
x"fbb00",-- -1104
x"01500",-- 336
x"fe400",-- -448
x"00c00",-- 192
x"01000",-- 256
x"fc000",-- -1024
x"07700",-- 1904
x"f8a00",-- -1888
x"04400",-- 1088
x"ff800",-- -128
x"ff900",-- -112
x"fff00",-- -16
x"ff000",-- -256
x"04000",-- 1024
x"f9c00",-- -1600
x"04a00",-- 1184
x"01200",-- 288
x"fc000",-- -1024
x"00c00",-- 192
x"01700",-- 368
x"ffb00",-- -80
x"00100",-- 16
x"00300",-- 48
x"02200",-- 544
x"fdf00",-- -528
x"00200",-- 32
x"ff900",-- -112
x"fe100",-- -496
x"01700",-- 368
x"00200",-- 32
x"03700",-- 880
x"fe300",-- -464
x"fdd00",-- -560
x"04900",-- 1168
x"fbb00",-- -1104
x"00700",-- 112
x"03e00",-- 992
x"fc000",-- -1024
x"03000",-- 768
x"fbf00",-- -1040
x"02b00",-- 688
x"fed00",-- -304
x"fcb00",-- -848
x"03600",-- 864
x"fef00",-- -272
x"fea00",-- -352
x"00800",-- 128
x"01c00",-- 448
x"fb200",-- -1248
x"02b00",-- 688
x"fd900",-- -624
x"ffd00",-- -48
x"ffb00",-- -80
x"ff200",-- -224
x"01f00",-- 496
x"fed00",-- -304
x"02000",-- 512
x"fd600",-- -672
x"fe400",-- -448
x"02d00",-- 720
x"fd700",-- -656
x"ff800",-- -128
x"04800",-- 1152
x"fc900",-- -880
x"02e00",-- 736
x"fed00",-- -304
x"fe100",-- -496
x"00600",-- 96
x"ffa00",-- -96
x"00e00",-- 224
x"fed00",-- -304
x"03e00",-- 992
x"fcd00",-- -816
x"02400",-- 576
x"ffc00",-- -64
x"fee00",-- -288
x"00d00",-- 208
x"00800",-- 128
x"00d00",-- 208
x"00000",-- 0
x"fec00",-- -320
x"01600",-- 352
x"fd700",-- -656
x"ffc00",-- -64
x"01500",-- 336
x"fc600",-- -928
x"04500",-- 1104
x"fff00",-- -16
x"00a00",-- 160
x"ffe00",-- -32
x"ff000",-- -256
x"ff400",-- -192
x"fe500",-- -432
x"01500",-- 336
x"00d00",-- 208
x"ff100",-- -240
x"00b00",-- 176
x"fe800",-- -384
x"01300",-- 304
x"ffb00",-- -80
x"fe200",-- -480
x"04400",-- 1088
x"fd800",-- -640
x"03c00",-- 960
x"ffa00",-- -96
x"feb00",-- -336
x"02a00",-- 672
x"fe200",-- -480
x"03e00",-- 992
x"ff100",-- -240
x"01f00",-- 496
x"00a00",-- 160
x"fe100",-- -496
x"02b00",-- 688
x"fd500",-- -688
x"01e00",-- 480
x"fc900",-- -880
x"01500",-- 336
x"01d00",-- 464
x"fc800",-- -896
x"04c00",-- 1216
x"fb400",-- -1216
x"01700",-- 368
x"fe600",-- -416
x"00d00",-- 208
x"ffe00",-- -32
x"fdc00",-- -576
x"02f00",-- 752
x"f9c00",-- -1600
x"04e00",-- 1248
x"fcf00",-- -784
x"ff200",-- -224
x"01000",-- 256
x"fc800",-- -896
x"02200",-- 544
x"fe800",-- -384
x"fef00",-- -272
x"01300",-- 304
x"fe700",-- -400
x"00500",-- 80
x"03000",-- 768
x"fc600",-- -928
x"03e00",-- 992
x"fd900",-- -624
x"fff00",-- -16
x"03300",-- 816
x"fe200",-- -480
x"02100",-- 528
x"ffd00",-- -48
x"00900",-- 144
x"00400",-- 64
x"02400",-- 576
x"00000",-- 0
x"00600",-- 96
x"00400",-- 64
x"01300",-- 304
x"01800",-- 384
x"fde00",-- -544
x"02f00",-- 752
x"ff500",-- -176
x"fef00",-- -272
x"03600",-- 864
x"fec00",-- -320
x"02300",-- 560
x"feb00",-- -336
x"ffe00",-- -32
x"02800",-- 640
x"fce00",-- -800
x"00200",-- 32
x"01200",-- 288
x"fc700",-- -912
x"00500",-- 80
x"00b00",-- 176
x"ff200",-- -224
x"00e00",-- 224
x"fe700",-- -400
x"00100",-- 16
x"fe800",-- -384
x"ffd00",-- -48
x"00100",-- 16
x"fe200",-- -480
x"00f00",-- 240
x"fed00",-- -304
x"01100",-- 272
x"fe700",-- -400
x"00600",-- 96
x"ff300",-- -208
x"01000",-- 256
x"ffb00",-- -80
x"ff200",-- -224
x"02d00",-- 720
x"fd200",-- -736
x"01000",-- 256
x"fe800",-- -384
x"ffd00",-- -48
x"00000",-- 0
x"ff900",-- -112
x"00f00",-- 240
x"fe400",-- -448
x"02300",-- 560
x"fe500",-- -432
x"fe800",-- -384
x"ff700",-- -144
x"fea00",-- -352
x"00800",-- 128
x"00800",-- 128
x"00a00",-- 160
x"00600",-- 96
x"fe600",-- -416
x"fdf00",-- -528
x"02a00",-- 672
x"feb00",-- -336
x"00100",-- 16
x"01000",-- 256
x"ff100",-- -240
x"00c00",-- 192
x"ffd00",-- -48
x"ff000",-- -256
x"ff300",-- -208
x"01100",-- 272
x"ff200",-- -224
x"02f00",-- 752
x"ffb00",-- -80
x"00100",-- 16
x"fff00",-- -16
x"fcf00",-- -784
x"02000",-- 512
x"ff400",-- -192
x"02100",-- 528
x"ff000",-- -256
x"fff00",-- -16
x"02800",-- 640
x"fda00",-- -608
x"01600",-- 352
x"fef00",-- -272
x"fea00",-- -352
x"03000",-- 768
x"00500",-- 80
x"01400",-- 320
x"00d00",-- 208
x"fe500",-- -432
x"fea00",-- -352
x"00b00",-- 176
x"00f00",-- 240
x"01700",-- 368
x"00600",-- 96
x"ffb00",-- -80
x"01900",-- 400
x"ff100",-- -240
x"fff00",-- -16
x"00900",-- 144
x"fec00",-- -320
x"01c00",-- 448
x"00c00",-- 192
x"00b00",-- 176
x"00300",-- 48
x"fdf00",-- -528
x"ffb00",-- -80
x"ffc00",-- -64
x"00800",-- 128
x"00800",-- 128
x"00100",-- 16
x"00300",-- 48
x"ffe00",-- -32
x"fef00",-- -272
x"ffb00",-- -80
x"ff200",-- -224
x"ffa00",-- -96
x"01000",-- 256
x"00e00",-- 224
x"00100",-- 16
x"ff100",-- -240
x"ff500",-- -176
x"ff000",-- -256
x"ffb00",-- -80
x"00300",-- 48
x"01500",-- 336
x"00500",-- 80
x"ff700",-- -144
x"ff900",-- -112
x"ff500",-- -176
x"ffc00",-- -64
x"ff700",-- -144
x"01e00",-- 480
x"00300",-- 48
x"01400",-- 320
x"01200",-- 288
x"fdb00",-- -592
x"00a00",-- 160
x"ffc00",-- -64
x"ffb00",-- -80
x"00100",-- 16
x"00a00",-- 160
x"00300",-- 48
x"ff400",-- -192
x"ffe00",-- -32
x"ff000",-- -256
x"fff00",-- -16
x"ffa00",-- -96
x"fff00",-- -16
x"01000",-- 256
x"00500",-- 80
x"fe500",-- -432
x"fe500",-- -432
x"fff00",-- -16
x"ff000",-- -256
x"00200",-- 32
x"00200",-- 32
x"00600",-- 96
x"01200",-- 288
x"00000",-- 0
x"fff00",-- -16
x"00200",-- 32
x"ffa00",-- -96
x"00900",-- 144
x"01b00",-- 432
x"00500",-- 80
x"01a00",-- 416
x"ffa00",-- -96
x"00200",-- 32
x"ffc00",-- -64
x"00e00",-- 224
x"01d00",-- 464
x"00200",-- 32
x"01900",-- 400
x"00a00",-- 160
x"00200",-- 32
x"ff500",-- -176
x"ffc00",-- -64
x"ff700",-- -144
x"ffe00",-- -32
x"00e00",-- 224
x"00c00",-- 192
x"00000",-- 0
x"fe600",-- -416
x"feb00",-- -336
x"ff600",-- -160
x"fff00",-- -16
x"00700",-- 112
x"ff300",-- -208
x"00000",-- 0
x"ff800",-- -128
x"ff200",-- -224
x"00000",-- 0
x"fe400",-- -448
x"00500",-- 80
x"00500",-- 80
x"00d00",-- 208
x"01600",-- 352
x"ff600",-- -160
x"ff200",-- -224
x"ffc00",-- -64
x"00200",-- 32
x"01200",-- 288
x"01600",-- 352
x"fe800",-- -384
x"ff900",-- -112
x"ff000",-- -256
x"ffa00",-- -96
x"00a00",-- 160
x"ff500",-- -176
x"ff900",-- -112
x"ff500",-- -176
x"ffd00",-- -48
x"00300",-- 48
x"ff200",-- -224
x"fe100",-- -496
x"ff100",-- -240
x"00300",-- 48
x"01300",-- 304
x"01300",-- 304
x"00100",-- 16
x"ff500",-- -176
x"ffd00",-- -48
x"01200",-- 288
x"01d00",-- 464
x"01f00",-- 496
x"01900",-- 400
x"00c00",-- 192
x"01600",-- 352
x"01700",-- 368
x"00d00",-- 208
x"01200",-- 288
x"00800",-- 128
x"00500",-- 80
x"01600",-- 352
x"00c00",-- 192
x"ff700",-- -144
x"fea00",-- -352
x"fec00",-- -320
x"ff800",-- -128
x"00500",-- 80
x"00300",-- 48
x"fe900",-- -368
x"fe100",-- -496
x"fe300",-- -464
x"feb00",-- -336
x"ff200",-- -224
x"fef00",-- -272
x"fe600",-- -416
x"ff400",-- -192
x"ff400",-- -192
x"ff500",-- -176
x"fef00",-- -272
x"fe700",-- -400
x"ff500",-- -176
x"00000",-- 0
x"00b00",-- 176
x"00900",-- 144
x"ffc00",-- -64
x"ff400",-- -192
x"ffd00",-- -48
x"00e00",-- 224
x"01600",-- 352
x"00f00",-- 240
x"00d00",-- 208
x"00b00",-- 176
x"00a00",-- 160
x"00e00",-- 224
x"00d00",-- 208
x"00800",-- 128
x"00c00",-- 192
x"01500",-- 336
x"01900",-- 400
x"01200",-- 288
x"00f00",-- 240
x"00500",-- 80
x"00900",-- 144
x"00f00",-- 240
x"01700",-- 368
x"00800",-- 128
x"00500",-- 80
x"fff00",-- -16
x"ff800",-- -128
x"00100",-- 16
x"ff900",-- -112
x"ffd00",-- -48
x"ffa00",-- -96
x"ff700",-- -144
x"ff900",-- -112
x"ff600",-- -160
x"fed00",-- -304
x"fed00",-- -304
x"fee00",-- -288
x"feb00",-- -336
x"ff300",-- -208
x"fed00",-- -304
x"fe300",-- -464
x"fe900",-- -368
x"fed00",-- -304
x"ff400",-- -192
x"ff300",-- -208
x"ff500",-- -176
x"ff100",-- -240
x"ff500",-- -176
x"ffa00",-- -96
x"ffe00",-- -32
x"00000",-- 0
x"00000",-- 0
x"00400",-- 64
x"00900",-- 144
x"00f00",-- 240
x"00e00",-- 224
x"01600",-- 352
x"01400",-- 320
x"01100",-- 272
x"00e00",-- 224
x"01700",-- 368
x"01a00",-- 416
x"01c00",-- 448
x"01d00",-- 464
x"01400",-- 320
x"01400",-- 320
x"00f00",-- 240
x"01200",-- 288
x"00f00",-- 240
x"00900",-- 144
x"00700",-- 112
x"fff00",-- -16
x"ffc00",-- -64
x"ff900",-- -112
x"ff100",-- -240
x"fee00",-- -288
x"fe700",-- -400
x"fe600",-- -416
x"fe500",-- -432
x"fe300",-- -464
x"fe300",-- -464
x"fe400",-- -448
x"fe300",-- -464
x"fe600",-- -416
x"fe700",-- -400
x"fe400",-- -448
x"fec00",-- -320
x"fee00",-- -288
x"ff400",-- -192
x"ff500",-- -176
x"ff800",-- -128
x"ff700",-- -144
x"ff900",-- -112
x"00400",-- 64
x"00400",-- 64
x"00d00",-- 208
x"00b00",-- 176
x"00f00",-- 240
x"00d00",-- 208
x"01000",-- 256
x"00e00",-- 224
x"01300",-- 304
x"01300",-- 304
x"01100",-- 272
x"01300",-- 304
x"00c00",-- 192
x"00d00",-- 208
x"00700",-- 112
x"00b00",-- 176
x"00800",-- 128
x"00800",-- 128
x"00400",-- 64
x"00100",-- 16
x"ffc00",-- -64
x"ff800",-- -128
x"ffa00",-- -96
x"ff500",-- -176
x"ff900",-- -112
x"ff400",-- -192
x"ff300",-- -208
x"ff200",-- -224
x"fed00",-- -304
x"ff000",-- -256
x"fee00",-- -288
x"fef00",-- -272
x"ff200",-- -224
x"ff500",-- -176
x"ff300",-- -208
x"ff500",-- -176
x"ff200",-- -224
x"ff700",-- -144
x"ffa00",-- -96
x"fff00",-- -16
x"fff00",-- -16
x"00200",-- 32
x"00400",-- 64
x"00100",-- 16
x"00600",-- 96
x"00700",-- 112
x"00b00",-- 176
x"00c00",-- 192
x"00e00",-- 224
x"00f00",-- 240
x"00e00",-- 224
x"00e00",-- 224
x"00f00",-- 240
x"00e00",-- 224
x"00f00",-- 240
x"00f00",-- 240
x"00b00",-- 176
x"00a00",-- 160
x"00800",-- 128
x"00500",-- 80
x"00400",-- 64
x"00300",-- 48
x"00100",-- 16
x"ffe00",-- -32
x"ffd00",-- -48
x"ffb00",-- -80
x"ff800",-- -128
x"ff600",-- -160
x"ff600",-- -160
x"ff500",-- -176
x"ff300",-- -208
x"ff400",-- -192
x"ff200",-- -224
x"ff300",-- -208
x"ff300",-- -208
x"ff300",-- -208
x"ff400",-- -192
x"ff500",-- -176
x"ff600",-- -160
x"ff700",-- -144
x"ff900",-- -112
x"ffb00",-- -80
x"ffd00",-- -48
x"ffd00",-- -48
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00300",-- 48
x"00700",-- 112
x"00600",-- 96
x"00800",-- 128
x"00600",-- 96
x"00700",-- 112
x"00600",-- 96
x"00900",-- 144
x"00900",-- 144
x"00700",-- 112
x"00a00",-- 160
x"00600",-- 96
x"00700",-- 112
x"00400",-- 64
x"00500",-- 80
x"00300",-- 48
x"00400",-- 64
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"ffd00",-- -48
x"ffd00",-- -48
x"ffc00",-- -64
x"ffe00",-- -32
x"ffc00",-- -64
x"ffb00",-- -80
x"ffa00",-- -96
x"ff900",-- -112
x"ff900",-- -112
x"ff900",-- -112
x"ffa00",-- -96
x"ff900",-- -112
x"ff900",-- -112
x"ffa00",-- -96
x"ffb00",-- -80
x"ffa00",-- -96
x"ffc00",-- -64
x"ff900",-- -112
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"00100",-- 16
x"00000",-- 0
x"00200",-- 32
x"00000",-- 0
x"00400",-- 64
x"00300",-- 48
x"00400",-- 64
x"00300",-- 48
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00200",-- 32
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00300",-- 48
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00200",-- 32
x"00000",-- 0
x"00200",-- 32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffd00",-- -48
x"ffe00",-- -32
x"ffc00",-- -64
x"fff00",-- -16
x"ffd00",-- -48
x"ffe00",-- -32
x"ffd00",-- -48
x"ffc00",-- -64
x"ffd00",-- -48
x"ffc00",-- -64
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00000",-- 0
x"00200",-- 32
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"00000",-- 0
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffd00",-- -48
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffd00",-- -48
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"00000",-- 0
x"ffe00",-- -32
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"ffe00",-- -32
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00200",-- 32
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00300",-- 48
x"00200",-- 32
x"00300",-- 48
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00300",-- 48
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"fff00",-- -16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"ffc00",-- -64
x"ffd00",-- -48
x"ff900",-- -112
x"ffa00",-- -96
x"ff500",-- -176
x"ff400",-- -192
x"fec00",-- -320
x"fea00",-- -352
x"fd200",-- -736
x"f9e00",-- -1568
x"fd000",-- -768
x"00700",-- 112
x"fef00",-- -272
x"fca00",-- -864
x"fa500",-- -1456
x"fae00",-- -1312
x"ff000",-- -256
x"00800",-- 128
x"ff000",-- -256
x"fc400",-- -960
x"fbb00",-- -1104
x"ffe00",-- -32
x"03a00",-- 928
x"03e00",-- 992
x"01900",-- 400
x"00800",-- 128
x"04100",-- 1040
x"08300",-- 2096
x"09300",-- 2352
x"07900",-- 1936
x"06b00",-- 1712
x"07e00",-- 2016
x"09600",-- 2400
x"09400",-- 2368
x"08300",-- 2096
x"06700",-- 1648
x"05400",-- 1344
x"05700",-- 1392
x"04200",-- 1056
x"02000",-- 512
x"01600",-- 352
x"01500",-- 336
x"ffb00",-- -80
x"fd700",-- -656
x"fcf00",-- -784
x"fce00",-- -800
x"fca00",-- -864
x"fcc00",-- -832
x"fb700",-- -1168
x"f9700",-- -1680
x"fa300",-- -1488
x"fc200",-- -992
x"fc300",-- -976
x"fb500",-- -1200
x"faa00",-- -1376
x"fa900",-- -1392
x"fbe00",-- -1056
x"fdb00",-- -592
x"fdb00",-- -592
x"fc600",-- -928
x"fc500",-- -944
x"fd500",-- -688
x"fe300",-- -464
x"fee00",-- -288
x"fed00",-- -304
x"fe400",-- -448
x"fe300",-- -464
x"ff100",-- -240
x"ffb00",-- -80
x"00000",-- 0
x"00400",-- 64
x"00200",-- 32
x"00000",-- 0
x"00500",-- 80
x"01200",-- 288
x"01c00",-- 448
x"01d00",-- 464
x"01700",-- 368
x"01400",-- 320
x"01700",-- 368
x"02100",-- 528
x"02a00",-- 672
x"02300",-- 560
x"01700",-- 368
x"01300",-- 304
x"01700",-- 368
x"01b00",-- 432
x"01e00",-- 480
x"01500",-- 336
x"00400",-- 64
x"00300",-- 48
x"00800",-- 128
x"00700",-- 112
x"00300",-- 48
x"ffc00",-- -64
x"ff100",-- -240
x"fec00",-- -320
x"ff300",-- -208
x"ff400",-- -192
x"fee00",-- -288
x"fed00",-- -304
x"fe900",-- -368
x"fe300",-- -464
x"fe900",-- -368
x"ff200",-- -224
x"fef00",-- -272
x"fed00",-- -304
x"fee00",-- -288
x"fec00",-- -320
x"ff100",-- -240
x"ffd00",-- -48
x"fff00",-- -16
x"ff900",-- -112
x"ffa00",-- -96
x"ffe00",-- -32
x"00300",-- 48
x"00a00",-- 160
x"00e00",-- 224
x"00700",-- 112
x"00400",-- 64
x"00a00",-- 160
x"00e00",-- 224
x"01000",-- 256
x"00f00",-- 240
x"00c00",-- 192
x"00800",-- 128
x"00900",-- 144
x"00e00",-- 224
x"00d00",-- 208
x"00a00",-- 160
x"00700",-- 112
x"00200",-- 32
x"00000",-- 0
x"00000",-- 0
x"00200",-- 32
x"ffe00",-- -32
x"ff700",-- -144
x"ff800",-- -128
x"ff400",-- -192
x"ff600",-- -160
x"ff900",-- -112
x"ff700",-- -144
x"ff300",-- -208
x"ff200",-- -224
x"ff400",-- -192
x"ff600",-- -160
x"ff600",-- -160
x"ff900",-- -112
x"ff500",-- -176
x"ff300",-- -208
x"ff700",-- -144
x"ffb00",-- -80
x"ff800",-- -128
x"fff00",-- -16
x"fec00",-- -320
x"fd400",-- -704
x"fef00",-- -272
x"00600",-- 96
x"ffa00",-- -96
x"fd800",-- -640
x"fc400",-- -960
x"fd200",-- -736
x"ff000",-- -256
x"fee00",-- -288
x"fce00",-- -800
x"fad00",-- -1328
x"fb600",-- -1184
x"fd700",-- -656
x"fe300",-- -464
x"fcf00",-- -784
x"fba00",-- -1120
x"fc200",-- -992
x"fdd00",-- -560
x"ff000",-- -256
x"ffc00",-- -64
x"00000",-- 0
x"00300",-- 48
x"02000",-- 512
x"03f00",-- 1008
x"04300",-- 1072
x"05700",-- 1392
x"07200",-- 1824
x"07500",-- 1872
x"06b00",-- 1712
x"07600",-- 1888
x"08f00",-- 2288
x"0b000",-- 2816
x"0c200",-- 3104
x"0a100",-- 2576
x"07700",-- 1904
x"08200",-- 2080
x"0ac00",-- 2752
x"0ac00",-- 2752
x"07b00",-- 1968
x"04400",-- 1088
x"02b00",-- 688
x"03100",-- 784
x"03d00",-- 976
x"02600",-- 608
x"fed00",-- -304
x"fbe00",-- -1056
x"fb700",-- -1168
x"fc500",-- -944
x"fc200",-- -992
x"fae00",-- -1312
x"f9b00",-- -1616
x"f8800",-- -1920
x"f8100",-- -2032
x"f9900",-- -1648
x"fac00",-- -1344
x"fa300",-- -1488
x"f9800",-- -1664
x"f9700",-- -1680
x"f9800",-- -1664
x"fa700",-- -1424
x"fca00",-- -864
x"fd100",-- -752
x"fba00",-- -1120
x"fb600",-- -1184
x"fc800",-- -896
x"fdb00",-- -592
x"ff200",-- -224
x"ff800",-- -128
x"fe400",-- -448
x"fd800",-- -640
x"fef00",-- -272
x"00d00",-- 208
x"01500",-- 336
x"00e00",-- 224
x"00500",-- 80
x"00200",-- 32
x"01100",-- 272
x"02900",-- 656
x"03100",-- 784
x"02100",-- 528
x"01600",-- 352
x"01c00",-- 448
x"02500",-- 592
x"02e00",-- 736
x"03200",-- 800
x"02800",-- 640
x"01300",-- 304
x"01100",-- 272
x"01e00",-- 480
x"02000",-- 512
x"01700",-- 368
x"00f00",-- 240
x"00000",-- 0
x"ff400",-- -192
x"00000",-- 0
x"00a00",-- 160
x"ffd00",-- -48
x"fe500",-- -432
x"fdc00",-- -576
x"fdf00",-- -528
x"fd700",-- -656
x"fdd00",-- -560
x"fdc00",-- -576
x"fc700",-- -912
x"fb800",-- -1152
x"fb900",-- -1136
x"fc400",-- -960
x"fc500",-- -944
x"fbd00",-- -1072
x"fad00",-- -1328
x"fa100",-- -1520
x"fa900",-- -1392
x"fb900",-- -1136
x"fbc00",-- -1088
x"fb600",-- -1184
x"fad00",-- -1328
x"fb500",-- -1200
x"fc700",-- -912
x"fd600",-- -672
x"fe200",-- -480
x"fea00",-- -352
x"ff600",-- -160
x"00900",-- 144
x"02d00",-- 720
x"04a00",-- 1184
x"05300",-- 1328
x"04500",-- 1104
x"07700",-- 1904
x"0b300",-- 2864
x"09d00",-- 2512
x"07d00",-- 2000
x"09500",-- 2384
x"0bd00",-- 3024
x"0cf00",-- 3312
x"0e700",-- 3696
x"0db00",-- 3504
x"09f00",-- 2544
x"08e00",-- 2272
x"0d300",-- 3376
x"0e400",-- 3648
x"09500",-- 2384
x"05700",-- 1392
x"05200",-- 1312
x"04400",-- 1088
x"02c00",-- 704
x"02f00",-- 752
x"00c00",-- 192
x"fb500",-- -1200
x"f9600",-- -1696
x"fba00",-- -1120
x"faf00",-- -1296
x"f8100",-- -2032
x"f8700",-- -1936
x"f7f00",-- -2064
x"f4d00",-- -2864
x"f5100",-- -2800
x"f8e00",-- -1824
x"f8c00",-- -1856
x"f6000",-- -2560
x"f6b00",-- -2384
x"f7a00",-- -2144
x"f7000",-- -2304
x"f9300",-- -1744
x"fc700",-- -912
x"fad00",-- -1328
x"f8500",-- -1968
x"fac00",-- -1344
x"fdd00",-- -560
x"fdc00",-- -576
x"fe300",-- -464
x"ff500",-- -176
x"fe000",-- -512
x"fd600",-- -672
x"01100",-- 272
x"03500",-- 848
x"01200",-- 288
x"00800",-- 128
x"02400",-- 576
x"02700",-- 624
x"02500",-- 592
x"04f00",-- 1264
x"05100",-- 1296
x"02400",-- 576
x"01e00",-- 480
x"04d00",-- 1232
x"04000",-- 1024
x"02900",-- 656
x"02500",-- 592
x"ffe00",-- -32
x"00500",-- 80
x"02300",-- 560
x"01400",-- 320
x"fd300",-- -720
x"fbb00",-- -1104
x"fc700",-- -912
x"fd300",-- -720
x"fbf00",-- -1040
x"f9700",-- -1680
x"f7c00",-- -2112
x"f7800",-- -2176
x"f8400",-- -1984
x"f8e00",-- -1824
x"f8e00",-- -1824
x"f7500",-- -2224
x"f7600",-- -2208
x"f9b00",-- -1616
x"fb200",-- -1248
x"fc500",-- -944
x"fe300",-- -464
x"ffb00",-- -80
x"00900",-- 144
x"03f00",-- 1008
x"06700",-- 1648
x"07d00",-- 2000
x"09400",-- 2368
x"0b400",-- 2880
x"0d500",-- 3408
x"0c900",-- 3216
x"0e400",-- 3648
x"12a00",-- 4768
x"14200",-- 5152
x"10c00",-- 4288
x"0dc00",-- 3520
x"0fc00",-- 4032
x"12400",-- 4672
x"0ff00",-- 4080
x"0c700",-- 3184
x"09900",-- 2448
x"06600",-- 1632
x"05800",-- 1408
x"06800",-- 1664
x"04200",-- 1056
x"fe100",-- -496
x"fad00",-- -1328
x"fbc00",-- -1088
x"fb100",-- -1264
x"f8d00",-- -1840
x"f8300",-- -2000
x"f7600",-- -2208
x"f4500",-- -2992
x"f3700",-- -3216
x"f6200",-- -2528
x"f6e00",-- -2336
x"f4900",-- -2928
x"f4200",-- -3040
x"f5300",-- -2768
x"f4a00",-- -2912
x"f5300",-- -2768
x"f8700",-- -1936
x"f9300",-- -1744
x"f6400",-- -2496
x"f6900",-- -2416
x"fa000",-- -1536
x"fae00",-- -1312
x"fae00",-- -1312
x"fc800",-- -896
x"fc300",-- -976
x"fa900",-- -1392
x"fcf00",-- -784
x"00e00",-- 224
x"00200",-- 32
x"fe300",-- -464
x"ffb00",-- -80
x"00a00",-- 160
x"01100",-- 272
x"01500",-- 336
x"02500",-- 592
x"03600",-- 864
x"01c00",-- 448
x"00700",-- 112
x"01200",-- 288
x"02800",-- 640
x"02d00",-- 720
x"01200",-- 288
x"fe600",-- -416
x"fdc00",-- -576
x"ff500",-- -176
x"00400",-- 64
x"fe400",-- -448
x"fb700",-- -1168
x"fb500",-- -1200
x"fc900",-- -880
x"fd400",-- -704
x"fdc00",-- -576
x"fd300",-- -720
x"fc800",-- -896
x"fe000",-- -512
x"00e00",-- 224
x"02200",-- 544
x"02900",-- 656
x"04100",-- 1040
x"06900",-- 1680
x"05300",-- 1328
x"05300",-- 1328
x"07c00",-- 1984
x"0c300",-- 3120
x"10300",-- 4144
x"0e200",-- 3616
x"0a100",-- 2576
x"0a300",-- 2608
x"0fa00",-- 4000
x"13a00",-- 5024
x"10700",-- 4208
x"09500",-- 2384
x"06800",-- 1664
x"08300",-- 2096
x"0ad00",-- 2768
x"09a00",-- 2464
x"04300",-- 1072
x"feb00",-- -336
x"fc700",-- -912
x"fe000",-- -512
x"fef00",-- -272
x"fd000",-- -768
x"f9b00",-- -1616
x"f7400",-- -2240
x"f6600",-- -2464
x"f7000",-- -2304
x"f9300",-- -1744
x"f9800",-- -1664
x"f7600",-- -2208
x"f5200",-- -2784
x"f5400",-- -2752
x"f7300",-- -2256
x"f9600",-- -1696
x"fa700",-- -1424
x"f8e00",-- -1824
x"f6d00",-- -2352
x"f7100",-- -2288
x"fa300",-- -1488
x"fcf00",-- -784
x"fc900",-- -880
x"fa500",-- -1456
x"f8c00",-- -1856
x"fa400",-- -1472
x"fd600",-- -672
x"ff800",-- -128
x"fe100",-- -496
x"fb900",-- -1136
x"f9d00",-- -1584
x"fde00",-- -544
x"fff00",-- -16
x"feb00",-- -336
x"ff100",-- -240
x"fd600",-- -672
x"fc200",-- -992
x"fd200",-- -736
x"fed00",-- -304
x"ff300",-- -208
x"ff300",-- -208
x"fca00",-- -864
x"fac00",-- -1344
x"fbd00",-- -1072
x"fed00",-- -304
x"ffd00",-- -48
x"fd800",-- -640
x"fb100",-- -1264
x"fae00",-- -1312
x"fe700",-- -400
x"01e00",-- 480
x"01900",-- 400
x"ff700",-- -144
x"fff00",-- -16
x"03100",-- 784
x"06600",-- 1632
x"08d00",-- 2256
x"09300",-- 2352
x"09c00",-- 2496
x"0ac00",-- 2752
x"0c100",-- 3088
x"09e00",-- 2528
x"0b900",-- 2960
x"14900",-- 5264
x"17500",-- 5968
x"0ea00",-- 3744
x"07e00",-- 2016
x"0dd00",-- 3536
x"16f00",-- 5872
x"15900",-- 5520
x"0c800",-- 3200
x"06b00",-- 1712
x"04d00",-- 1232
x"07100",-- 1808
x"0ad00",-- 2768
x"08300",-- 2096
x"fe100",-- -496
x"f6b00",-- -2384
x"f9500",-- -1712
x"fd400",-- -704
x"fab00",-- -1360
x"f7000",-- -2304
x"f5700",-- -2704
x"f2300",-- -3536
x"f0500",-- -4016
x"f4a00",-- -2912
x"f8c00",-- -1856
x"f5a00",-- -2656
x"f1000",-- -3840
x"f1b00",-- -3664
x"f4200",-- -3040
x"f5800",-- -2688
x"f8700",-- -1936
x"f9f00",-- -1552
x"f6300",-- -2512
x"f2400",-- -3520
x"f4000",-- -3072
x"fc800",-- -896
x"01500",-- 336
x"fbf00",-- -1040
x"f4100",-- -3056
x"f3e00",-- -3104
x"fc000",-- -1024
x"02b00",-- 688
x"fff00",-- -16
x"f9600",-- -1696
x"f6200",-- -2528
x"f9f00",-- -1552
x"01100",-- 272
x"01a00",-- 416
x"fce00",-- -800
x"fad00",-- -1328
x"fa900",-- -1392
x"fce00",-- -800
x"00300",-- 48
x"00500",-- 80
x"fe500",-- -432
x"fc800",-- -896
x"fcc00",-- -832
x"fe900",-- -368
x"01c00",-- 448
x"03000",-- 768
x"00d00",-- 208
x"ffa00",-- -96
x"01d00",-- 464
x"06500",-- 1616
x"08d00",-- 2256
x"09300",-- 2352
x"08c00",-- 2240
x"0b000",-- 2816
x"0db00",-- 3504
x"0eb00",-- 3760
x"0e100",-- 3600
x"0de00",-- 3552
x"14b00",-- 5296
x"18900",-- 6288
x"14400",-- 5184
x"0ef00",-- 3824
x"11800",-- 4480
x"17800",-- 6016
x"18100",-- 6160
x"10f00",-- 4336
x"0ba00",-- 2976
x"09b00",-- 2480
x"0a300",-- 2608
x"0b600",-- 2912
x"07200",-- 1824
x"00200",-- 32
x"faf00",-- -1296
x"f9d00",-- -1584
x"fa800",-- -1408
x"f8e00",-- -1824
x"f5100",-- -2800
x"f2000",-- -3584
x"f0f00",-- -3856
x"efe00",-- -4128
x"f0200",-- -4064
x"f1e00",-- -3616
x"f1d00",-- -3632
x"ef300",-- -4304
x"ef000",-- -4352
x"f0e00",-- -3872
x"f2500",-- -3504
x"f3e00",-- -3104
x"f5400",-- -2752
x"f4800",-- -2944
x"f2700",-- -3472
x"f5300",-- -2768
x"f9b00",-- -1616
x"f9a00",-- -1632
x"f7700",-- -2192
x"f7a00",-- -2144
x"f8b00",-- -1872
x"f9b00",-- -1616
x"fae00",-- -1312
x"fb900",-- -1136
x"faa00",-- -1376
x"f9e00",-- -1568
x"f9f00",-- -1552
x"fbd00",-- -1072
x"fc800",-- -896
x"fb900",-- -1136
x"fc100",-- -1008
x"fc700",-- -912
x"fc600",-- -928
x"fd400",-- -704
x"fe100",-- -496
x"fed00",-- -304
x"ff400",-- -192
x"ff800",-- -128
x"00400",-- 64
x"01200",-- 288
x"02d00",-- 720
x"05400",-- 1344
x"05800",-- 1408
x"06000",-- 1536
x"08000",-- 2048
x"0b300",-- 2864
x"0cd00",-- 3280
x"10300",-- 4144
x"10100",-- 4112
x"0d200",-- 3360
x"0df00",-- 3568
x"11f00",-- 4592
x"1a300",-- 6704
x"1af00",-- 6896
x"13400",-- 4928
x"0f400",-- 3904
x"15000",-- 5376
x"1b200",-- 6944
x"1ad00",-- 6864
x"12b00",-- 4784
x"0c100",-- 3088
x"0ab00",-- 2736
x"0c700",-- 3184
x"0d400",-- 3392
x"08c00",-- 2240
x"00b00",-- 176
x"faa00",-- -1376
x"f9200",-- -1760
x"f9c00",-- -1600
x"f8a00",-- -1888
x"f5800",-- -2688
x"f1100",-- -3824
x"ede00",-- -4640
x"ec800",-- -4992
x"ee800",-- -4480
x"f1800",-- -3712
x"f0300",-- -4048
x"ec100",-- -5104
x"ead00",-- -5424
x"ed000",-- -4864
x"f0800",-- -3968
x"f2f00",-- -3344
x"f0e00",-- -3872
x"ef400",-- -4288
x"ef700",-- -4240
x"f3500",-- -3248
x"f7900",-- -2160
x"f6d00",-- -2352
x"f4e00",-- -2848
x"f4d00",-- -2864
x"f5f00",-- -2576
x"f9700",-- -1680
x"fb500",-- -1200
x"f9700",-- -1680
x"f8200",-- -2016
x"f8200",-- -2016
x"fa600",-- -1440
x"fd600",-- -672
x"fd600",-- -672
x"fbc00",-- -1088
x"fb100",-- -1264
x"fcb00",-- -848
x"ff600",-- -160
x"01000",-- 256
x"00a00",-- 160
x"ff600",-- -160
x"00300",-- 48
x"03400",-- 832
x"06200",-- 1568
x"07400",-- 1856
x"06500",-- 1616
x"07000",-- 1792
x"0a400",-- 2624
x"0e200",-- 3616
x"10700",-- 4208
x"12400",-- 4672
x"11d00",-- 4560
x"0fb00",-- 4016
x"0f900",-- 3984
x"14d00",-- 5328
x"1e500",-- 7760
x"1dc00",-- 7616
x"14200",-- 5152
x"10200",-- 4128
x"16c00",-- 5824
x"1e600",-- 7776
x"1ca00",-- 7328
x"13100",-- 4880
x"0c300",-- 3120
x"0a300",-- 2608
x"0c000",-- 3072
x"0e500",-- 3664
x"09d00",-- 2512
x"ff200",-- -224
x"f7700",-- -2192
x"f7400",-- -2240
x"f9600",-- -1696
x"f8200",-- -2016
x"f4500",-- -2992
x"ee900",-- -4464
x"ea400",-- -5568
x"ea600",-- -5536
x"ee900",-- -4464
x"f1900",-- -3696
x"ee100",-- -4592
x"e8d00",-- -5936
x"e8b00",-- -5968
x"ec600",-- -5024
x"f0900",-- -3952
x"f0a00",-- -3936
x"eff00",-- -4112
x"edc00",-- -4672
x"ec600",-- -5024
x"f2900",-- -3440
x"f7e00",-- -2080
x"f6300",-- -2512
x"f2700",-- -3472
x"f2200",-- -3552
x"f5200",-- -2784
x"f9d00",-- -1584
x"fab00",-- -1360
x"f7900",-- -2160
x"f5700",-- -2704
x"f7d00",-- -2096
x"fb800",-- -1152
x"fdd00",-- -560
x"fd200",-- -736
x"fa800",-- -1408
x"fb500",-- -1200
x"fee00",-- -288
x"01c00",-- 448
x"02500",-- 592
x"01a00",-- 416
x"01600",-- 352
x"02f00",-- 752
x"05f00",-- 1520
x"09900",-- 2448
x"09900",-- 2448
x"08800",-- 2176
x"0a600",-- 2656
x"0d700",-- 3440
x"10800",-- 4224
x"14200",-- 5152
x"14f00",-- 5360
x"10d00",-- 4304
x"0e400",-- 3648
x"12b00",-- 4784
x"1ed00",-- 7888
x"21e00",-- 8672
x"16f00",-- 5872
x"0f400",-- 3904
x"15c00",-- 5568
x"1f000",-- 7936
x"1fa00",-- 8096
x"16800",-- 5760
x"0e000",-- 3584
x"0ad00",-- 2768
x"0c100",-- 3088
x"0ea00",-- 3744
x"0c200",-- 3104
x"03100",-- 784
x"f9200",-- -1760
x"f6600",-- -2464
x"f8b00",-- -1872
x"f8700",-- -1936
x"f5500",-- -2736
x"f0500",-- -4016
x"ea600",-- -5536
x"e8200",-- -6112
x"ebb00",-- -5200
x"f0f00",-- -3856
x"ee900",-- -4464
x"e8800",-- -6016
x"e6400",-- -6592
x"e9700",-- -5776
x"ecf00",-- -4880
x"ef300",-- -4304
x"eea00",-- -4448
x"ebb00",-- -5200
x"ec100",-- -5104
x"ef200",-- -4320
x"f2500",-- -3504
x"f4a00",-- -2912
x"f3f00",-- -3088
x"f1a00",-- -3680
x"f2100",-- -3568
x"f4c00",-- -2880
x"f7400",-- -2240
x"f9400",-- -1728
x"f8500",-- -1968
x"f6000",-- -2560
x"f7300",-- -2256
x"fc500",-- -944
x"fed00",-- -304
x"fe200",-- -480
x"fcb00",-- -848
x"fd400",-- -704
x"00e00",-- 224
x"04200",-- 1056
x"05900",-- 1424
x"04300",-- 1072
x"04000",-- 1024
x"07100",-- 1808
x"0a200",-- 2592
x"0b600",-- 2912
x"0c600",-- 3168
x"0d200",-- 3360
x"0ed00",-- 3792
x"10600",-- 4192
x"14c00",-- 5312
x"15800",-- 5504
x"13e00",-- 5088
x"11a00",-- 4512
x"14100",-- 5136
x"1d800",-- 7552
x"20600",-- 8288
x"19700",-- 6512
x"13c00",-- 5056
x"17900",-- 6032
x"1dc00",-- 7616
x"1e500",-- 7760
x"16300",-- 5680
x"10000",-- 4096
x"0d500",-- 3408
x"0c700",-- 3184
x"0cf00",-- 3312
x"09e00",-- 2528
x"02300",-- 560
x"fa400",-- -1472
x"f7900",-- -2160
x"f7600",-- -2208
x"f5c00",-- -2624
x"f3500",-- -3248
x"ef000",-- -4352
x"eab00",-- -5456
x"e8a00",-- -5984
x"ea700",-- -5520
x"ed400",-- -4800
x"ec500",-- -5040
x"e8200",-- -6112
x"e7100",-- -6384
x"e7f00",-- -6160
x"ea100",-- -5616
x"ecc00",-- -4928
x"ee100",-- -4592
x"ed900",-- -4720
x"eb800",-- -5248
x"eb300",-- -5328
x"f0100",-- -4080
x"f5c00",-- -2624
x"f4100",-- -3056
x"f0400",-- -4032
x"eec00",-- -4416
x"f2200",-- -3552
x"f8900",-- -1904
x"fa800",-- -1408
x"f6500",-- -2480
x"f4000",-- -3072
x"f7000",-- -2304
x"fcb00",-- -848
x"00200",-- 32
x"fe900",-- -368
x"fbe00",-- -1056
x"fe100",-- -496
x"02900",-- 656
x"06100",-- 1552
x"06b00",-- 1712
x"05a00",-- 1440
x"05900",-- 1424
x"09100",-- 2320
x"0bc00",-- 3008
x"0dd00",-- 3536
x"0e800",-- 3712
x"0ec00",-- 3776
x"0ff00",-- 4080
x"12e00",-- 4832
x"16d00",-- 5840
x"15e00",-- 5600
x"13400",-- 4928
x"11c00",-- 4544
x"19000",-- 6400
x"21500",-- 8528
x"1de00",-- 7648
x"15c00",-- 5568
x"14f00",-- 5360
x"1c100",-- 7184
x"1e400",-- 7744
x"16400",-- 5696
x"15d00",-- 5584
x"15700",-- 5488
x"0b600",-- 2912
x"06d00",-- 1744
x"0a700",-- 2672
x"0ab00",-- 2736
x"02b00",-- 688
x"f7300",-- -2256
x"f4100",-- -3056
x"f4800",-- -2944
x"f5500",-- -2736
x"f4500",-- -2992
x"ee300",-- -4560
x"e8200",-- -6112
x"e5b00",-- -6736
x"eb100",-- -5360
x"eef00",-- -4368
x"ebf00",-- -5136
x"e7700",-- -6288
x"e4b00",-- -6992
x"e7600",-- -6304
x"ebf00",-- -5136
x"f0200",-- -4064
x"ef800",-- -4224
x"ea000",-- -5632
x"e8800",-- -6016
x"edc00",-- -4672
x"f5500",-- -2736
x"f7100",-- -2288
x"f0300",-- -4048
x"eb200",-- -5344
x"f0f00",-- -3856
x"f8100",-- -2032
x"f9d00",-- -1584
x"f7900",-- -2160
x"f4600",-- -2976
x"f3600",-- -3232
x"fa300",-- -1488
x"01500",-- 336
x"ff700",-- -144
x"fbf00",-- -1040
x"fcb00",-- -848
x"00800",-- 128
x"05000",-- 1280
x"07c00",-- 1984
x"07300",-- 1840
x"04500",-- 1104
x"06300",-- 1584
x"0bc00",-- 3008
x"0e000",-- 3584
x"0e800",-- 3712
x"0e200",-- 3616
x"0f400",-- 3904
x"10d00",-- 4304
x"16800",-- 5760
x"17e00",-- 6112
x"14100",-- 5136
x"12100",-- 4624
x"14700",-- 5232
x"1dc00",-- 7616
x"21700",-- 8560
x"19e00",-- 6624
x"14600",-- 5216
x"17d00",-- 6096
x"1d400",-- 7488
x"1f200",-- 7968
x"17500",-- 5968
x"0fe00",-- 4064
x"0d200",-- 3360
x"0d800",-- 3456
x"0d300",-- 3376
x"08500",-- 2128
x"02500",-- 592
x"fb300",-- -1232
x"f7300",-- -2256
x"f7000",-- -2304
x"f4c00",-- -2880
x"f2600",-- -3488
x"edf00",-- -4624
x"ea200",-- -5600
x"e8500",-- -6064
x"e9200",-- -5856
x"ebc00",-- -5184
x"eb000",-- -5376
x"e6d00",-- -6448
x"e4100",-- -7152
x"e6400",-- -6592
x"ebc00",-- -5184
x"eeb00",-- -4432
x"eb400",-- -5312
x"e7f00",-- -6160
x"ea000",-- -5632
x"ef700",-- -4240
x"f3200",-- -3296
x"f3100",-- -3312
x"edf00",-- -4624
x"ece00",-- -4896
x"f2800",-- -3456
x"f7700",-- -2192
x"f7700",-- -2192
x"f5200",-- -2784
x"f3700",-- -3216
x"f6000",-- -2560
x"fbc00",-- -1088
x"ff100",-- -240
x"fda00",-- -608
x"fc100",-- -1008
x"fdb00",-- -592
x"02100",-- 528
x"06000",-- 1536
x"06f00",-- 1776
x"05800",-- 1408
x"05800",-- 1408
x"08900",-- 2192
x"0ce00",-- 3296
x"0dc00",-- 3520
x"0db00",-- 3504
x"0e400",-- 3648
x"10700",-- 4208
x"12e00",-- 4832
x"16300",-- 5680
x"16f00",-- 5872
x"14a00",-- 5280
x"12a00",-- 4768
x"14500",-- 5200
x"1cb00",-- 7344
x"21600",-- 8544
x"1b200",-- 6944
x"14000",-- 5120
x"16b00",-- 5808
x"1ca00",-- 7328
x"20100",-- 8208
x"18e00",-- 6368
x"10300",-- 4144
x"0cd00",-- 3280
x"0d000",-- 3328
x"0de00",-- 3552
x"0a500",-- 2640
x"03000",-- 768
x"fb800",-- -1152
x"f7200",-- -2272
x"f7200",-- -2272
x"f5f00",-- -2576
x"f3900",-- -3184
x"eea00",-- -4448
x"e9200",-- -5856
x"e8000",-- -6144
x"e9f00",-- -5648
x"ec500",-- -5040
x"eb400",-- -5312
x"e6100",-- -6640
x"e2300",-- -7632
x"e5b00",-- -6736
x"edb00",-- -4688
x"ef900",-- -4208
x"e9500",-- -5808
x"e5d00",-- -6704
x"e9400",-- -5824
x"f1600",-- -3744
x"f4500",-- -2992
x"f1100",-- -3824
x"ec000",-- -5120
x"ec200",-- -5088
x"f3a00",-- -3168
x"f8a00",-- -1888
x"f7200",-- -2272
x"f3b00",-- -3152
x"f2f00",-- -3344
x"f6a00",-- -2400
x"fc900",-- -880
x"ffc00",-- -64
x"fd700",-- -656
x"fb800",-- -1152
x"fe000",-- -512
x"02c00",-- 704
x"07100",-- 1808
x"07900",-- 1936
x"05200",-- 1312
x"05400",-- 1344
x"09300",-- 2352
x"0d500",-- 3408
x"0eb00",-- 3760
x"0dc00",-- 3520
x"0df00",-- 3568
x"11200",-- 4384
x"13400",-- 4928
x"16200",-- 5664
x"16a00",-- 5792
x"14b00",-- 5296
x"12700",-- 4720
x"15100",-- 5392
x"1c700",-- 7280
x"20c00",-- 8384
x"1ad00",-- 6864
x"14500",-- 5200
x"16f00",-- 5872
x"1c700",-- 7280
x"1f200",-- 7968
x"18300",-- 6192
x"10100",-- 4112
x"0cb00",-- 3248
x"0cf00",-- 3312
x"0d900",-- 3472
x"09a00",-- 2464
x"02300",-- 560
x"fb400",-- -1216
x"f7600",-- -2208
x"f7100",-- -2288
x"f5a00",-- -2656
x"f2c00",-- -3392
x"ee600",-- -4512
x"e9300",-- -5840
x"e7e00",-- -6176
x"e9f00",-- -5648
x"ebd00",-- -5168
x"ea400",-- -5568
x"e2b00",-- -7504
x"e3000",-- -7424
x"ebc00",-- -5184
x"ed100",-- -4848
x"e9300",-- -5840
x"e7900",-- -6256
x"e7900",-- -6256
x"ecd00",-- -4912
x"f3300",-- -3280
x"efd00",-- -4144
x"eb500",-- -5296
x"ed300",-- -4816
x"f1d00",-- -3632
x"f5700",-- -2704
x"f6600",-- -2464
x"f4500",-- -2992
x"f2b00",-- -3408
x"f6300",-- -2512
x"fb800",-- -1152
x"fd600",-- -672
x"fce00",-- -800
x"fcb00",-- -848
x"fe600",-- -416
x"00c00",-- 192
x"04a00",-- 1184
x"07700",-- 1904
x"05200",-- 1312
x"04600",-- 1120
x"08700",-- 2160
x"0c000",-- 3072
x"0c600",-- 3168
x"0d200",-- 3360
x"0d300",-- 3376
x"0f200",-- 3872
x"13000",-- 4864
x"14a00",-- 5280
x"15500",-- 5456
x"12f00",-- 4848
x"13500",-- 4944
x"15000",-- 5376
x"17b00",-- 6064
x"1bd00",-- 7120
x"1d100",-- 7440
x"17700",-- 6000
x"14e00",-- 5344
x"19700",-- 6512
x"1db00",-- 7600
x"1b600",-- 7008
x"14000",-- 5120
x"0ef00",-- 3824
x"0cc00",-- 3264
x"0dc00",-- 3520
x"0d300",-- 3376
x"06700",-- 1648
x"fe800",-- -384
x"fa100",-- -1520
x"f8500",-- -1968
x"f7900",-- -2160
x"f5500",-- -2736
x"f0d00",-- -3888
x"eba00",-- -5216
x"e9700",-- -5776
x"ea000",-- -5632
x"ebc00",-- -5184
x"ea900",-- -5488
x"e5500",-- -6832
x"e3d00",-- -7216
x"e9c00",-- -5696
x"ec300",-- -5072
x"e9900",-- -5744
x"e7d00",-- -6192
x"e8600",-- -6048
x"ec400",-- -5056
x"f0600",-- -4000
x"ef500",-- -4272
x"ec300",-- -5072
x"ee400",-- -4544
x"f1f00",-- -3600
x"f2800",-- -3456
x"f4800",-- -2944
x"f5900",-- -2672
x"f4500",-- -2992
x"f5e00",-- -2592
x"f9400",-- -1728
x"fb300",-- -1232
x"fce00",-- -800
x"fe300",-- -464
x"fe700",-- -400
x"ff500",-- -176
x"02700",-- 624
x"05f00",-- 1520
x"05e00",-- 1504
x"05600",-- 1376
x"06c00",-- 1728
x"09c00",-- 2496
x"0bc00",-- 3008
x"0c200",-- 3104
x"0d900",-- 3472
x"0e800",-- 3712
x"10b00",-- 4272
x"12900",-- 4752
x"14e00",-- 5344
x"14700",-- 5232
x"12600",-- 4704
x"14200",-- 5152
x"15f00",-- 5616
x"18e00",-- 6368
x"1c300",-- 7216
x"19a00",-- 6560
x"15e00",-- 5600
x"17500",-- 5968
x"1ad00",-- 6864
x"1c200",-- 7200
x"17800",-- 6016
x"12000",-- 4608
x"0e100",-- 3600
x"0d500",-- 3408
x"0e300",-- 3632
x"0a200",-- 2592
x"02c00",-- 704
x"fd000",-- -768
x"f9f00",-- -1552
x"f8e00",-- -1824
x"f6f00",-- -2320
x"f3f00",-- -3088
x"ee700",-- -4496
x"eb300",-- -5328
x"ead00",-- -5424
x"ebb00",-- -5200
x"eb700",-- -5264
x"e7100",-- -6384
x"e6300",-- -6608
x"e9800",-- -5760
x"ea800",-- -5504
x"e9300",-- -5840
x"e9100",-- -5872
x"e9900",-- -5744
x"eba00",-- -5216
x"ee300",-- -4560
x"ee300",-- -4560
x"ecb00",-- -4944
x"ee900",-- -4464
x"f1200",-- -3808
x"f1d00",-- -3632
x"f3000",-- -3328
x"f4400",-- -3008
x"f4400",-- -3008
x"f5a00",-- -2656
x"f8100",-- -2032
x"fa000",-- -1536
x"fb400",-- -1216
x"fce00",-- -800
x"fe100",-- -496
x"ff400",-- -192
x"01a00",-- 416
x"04100",-- 1040
x"04b00",-- 1200
x"05400",-- 1344
x"07400",-- 1856
x"08e00",-- 2272
x"0ab00",-- 2736
x"0b700",-- 2928
x"0c900",-- 3216
x"0e800",-- 3712
x"10d00",-- 4304
x"11f00",-- 4592
x"12700",-- 4720
x"14000",-- 5120
x"14400",-- 5184
x"14400",-- 5184
x"14e00",-- 5344
x"16b00",-- 5808
x"1a600",-- 6752
x"1b600",-- 7008
x"17800",-- 6016
x"16200",-- 5664
x"18c00",-- 6336
x"1b600",-- 7008
x"19700",-- 6512
x"13600",-- 4960
x"0f400",-- 3904
x"0de00",-- 3552
x"0da00",-- 3488
x"0b700",-- 2928
x"05300",-- 1328
x"feb00",-- -336
x"fad00",-- -1328
x"f9d00",-- -1584
x"f8200",-- -2016
x"f3f00",-- -3088
x"efe00",-- -4128
x"ecd00",-- -4912
x"ebd00",-- -5168
x"eb800",-- -5248
x"ead00",-- -5424
x"e8700",-- -6032
x"e7500",-- -6320
x"e8700",-- -6032
x"e9d00",-- -5680
x"ea200",-- -5600
x"e8e00",-- -5920
x"e9500",-- -5808
x"eb400",-- -5312
x"ec800",-- -4992
x"ee400",-- -4544
x"ee300",-- -4560
x"ed200",-- -4832
x"efe00",-- -4128
x"f2200",-- -3552
x"f2200",-- -3552
x"f3d00",-- -3120
x"f4d00",-- -2864
x"f4700",-- -2960
x"f6c00",-- -2368
x"fa000",-- -1536
x"fad00",-- -1328
x"fc200",-- -992
x"fde00",-- -544
x"fed00",-- -304
x"01000",-- 256
x"03200",-- 800
x"04800",-- 1152
x"05a00",-- 1440
x"06800",-- 1664
x"07e00",-- 2016
x"0a200",-- 2592
x"0b700",-- 2928
x"0bb00",-- 2992
x"0d500",-- 3408
x"0f600",-- 3936
x"11200",-- 4384
x"12400",-- 4672
x"14200",-- 5152
x"13600",-- 4960
x"12600",-- 4704
x"13d00",-- 5072
x"16200",-- 5664
x"19900",-- 6544
x"1ac00",-- 6848
x"16c00",-- 5824
x"14500",-- 5200
x"17e00",-- 6112
x"1bc00",-- 7104
x"1a300",-- 6704
x"13d00",-- 5072
x"0f300",-- 3888
x"0df00",-- 3568
x"0e800",-- 3712
x"0cd00",-- 3280
x"07400",-- 1856
x"ffc00",-- -64
x"fbb00",-- -1104
x"fad00",-- -1328
x"f9600",-- -1696
x"f5800",-- -2688
x"f1900",-- -3696
x"edc00",-- -4672
x"ebe00",-- -5152
x"ec100",-- -5104
x"ebd00",-- -5168
x"ea700",-- -5520
x"e8700",-- -6032
x"e8200",-- -6112
x"e8500",-- -6064
x"ea800",-- -5504
x"eb800",-- -5248
x"ea400",-- -5568
x"e9e00",-- -5664
x"ebe00",-- -5152
x"ed700",-- -4752
x"ef600",-- -4256
x"f0100",-- -4080
x"eed00",-- -4400
x"efd00",-- -4144
x"f2300",-- -3536
x"f4400",-- -3008
x"f5600",-- -2720
x"f5500",-- -2736
x"f5a00",-- -2656
x"f7a00",-- -2144
x"fa800",-- -1408
x"fcc00",-- -832
x"fdd00",-- -560
x"fe000",-- -512
x"ff300",-- -208
x"02000",-- 512
x"04800",-- 1152
x"05700",-- 1392
x"06000",-- 1536
x"06900",-- 1680
x"08400",-- 2112
x"0ae00",-- 2784
x"0c500",-- 3152
x"0cf00",-- 3312
x"0d400",-- 3392
x"10100",-- 4112
x"11800",-- 4480
x"13800",-- 4992
x"14000",-- 5120
x"11800",-- 4480
x"12c00",-- 4800
x"16700",-- 5744
x"17700",-- 6000
x"19400",-- 6464
x"18600",-- 6240
x"16000",-- 5632
x"17000",-- 5888
x"19100",-- 6416
x"1a100",-- 6672
x"16500",-- 5712
x"11900",-- 4496
x"0e600",-- 3680
x"0d900",-- 3472
x"0d400",-- 3392
x"09100",-- 2320
x"02d00",-- 720
x"fda00",-- -608
x"fa900",-- -1392
x"fa500",-- -1456
x"f7300",-- -2256
x"f3000",-- -3328
x"efb00",-- -4176
x"ecf00",-- -4880
x"ec700",-- -5008
x"eca00",-- -4960
x"eb100",-- -5360
x"e9500",-- -5808
x"e9500",-- -5808
x"e8f00",-- -5904
x"e8a00",-- -5984
x"eb500",-- -5296
x"ec900",-- -4976
x"ea600",-- -5536
x"ea200",-- -5600
x"ed100",-- -4848
x"ef000",-- -4352
x"ef500",-- -4272
x"f0600",-- -4000
x"ef500",-- -4272
x"f0200",-- -4064
x"f4300",-- -3024
x"f5700",-- -2704
x"f4600",-- -2976
x"f5100",-- -2800
x"f7900",-- -2160
x"f9400",-- -1728
x"fb600",-- -1184
x"fd300",-- -720
x"fd900",-- -624
x"fee00",-- -288
x"01100",-- 272
x"03700",-- 880
x"05400",-- 1344
x"05d00",-- 1488
x"06100",-- 1552
x"07800",-- 1920
x"0a500",-- 2640
x"0ce00",-- 3296
x"0cc00",-- 3264
x"0c700",-- 3184
x"0f300",-- 3888
x"11d00",-- 4560
x"13800",-- 4992
x"12c00",-- 4800
x"11100",-- 4368
x"13600",-- 4960
x"16400",-- 5696
x"16c00",-- 5824
x"18400",-- 6208
x"17900",-- 6032
x"16500",-- 5712
x"17d00",-- 6096
x"18900",-- 6288
x"18900",-- 6288
x"16400",-- 5696
x"13000",-- 4864
x"0fb00",-- 4016
x"0db00",-- 3504
x"0d000",-- 3328
x"09b00",-- 2480
x"04400",-- 1088
x"ff000",-- -256
x"fb400",-- -1216
x"fa400",-- -1472
x"f8800",-- -1920
x"f4200",-- -3040
x"f0300",-- -4048
x"edc00",-- -4672
x"ed100",-- -4848
x"ed500",-- -4784
x"ebe00",-- -5152
x"e9b00",-- -5712
x"e8e00",-- -5920
x"e9a00",-- -5728
x"e9e00",-- -5664
x"ead00",-- -5424
x"ebb00",-- -5200
x"eb000",-- -5376
x"ea300",-- -5584
x"ec400",-- -5056
x"ef800",-- -4224
x"efa00",-- -4192
x"efa00",-- -4192
x"efb00",-- -4176
x"f0000",-- -4096
x"f3900",-- -3184
x"f5e00",-- -2592
x"f4e00",-- -2848
x"f4b00",-- -2896
x"f6900",-- -2416
x"f9700",-- -1680
x"fbd00",-- -1072
x"fd200",-- -736
x"fd700",-- -656
x"fe300",-- -464
x"01300",-- 304
x"03d00",-- 976
x"04b00",-- 1200
x"05500",-- 1360
x"06900",-- 1680
x"08400",-- 2112
x"09a00",-- 2464
x"0bb00",-- 2992
x"0d000",-- 3328
x"0da00",-- 3488
x"0ec00",-- 3776
x"10600",-- 4192
x"13800",-- 4992
x"13700",-- 4976
x"10800",-- 4224
x"12700",-- 4720
x"16600",-- 5728
x"16c00",-- 5824
x"17900",-- 6032
x"17300",-- 5936
x"15900",-- 5520
x"17600",-- 5984
x"19100",-- 6416
x"18900",-- 6288
x"15a00",-- 5536
x"11d00",-- 4560
x"0f600",-- 3936
x"0ed00",-- 3792
x"0d400",-- 3392
x"08d00",-- 2256
x"03c00",-- 960
x"ffb00",-- -80
x"fc200",-- -992
x"fa900",-- -1392
x"f8900",-- -1904
x"f4b00",-- -2896
x"f1100",-- -3824
x"ee100",-- -4592
x"edf00",-- -4624
x"ee100",-- -4592
x"ec100",-- -5104
x"ea500",-- -5552
x"eac00",-- -5440
x"e8c00",-- -5952
x"e8b00",-- -5968
x"ed600",-- -4768
x"ece00",-- -4896
x"ea600",-- -5536
x"ebb00",-- -5200
x"eac00",-- -5440
x"ee000",-- -4608
x"f3a00",-- -3168
x"f1100",-- -3824
x"ed000",-- -4864
x"ef900",-- -4208
x"f3e00",-- -3104
x"f6200",-- -2528
x"f7300",-- -2256
x"f4d00",-- -2864
x"f4100",-- -3056
x"f9000",-- -1792
x"fd100",-- -752
x"fe300",-- -464
x"fdd00",-- -560
x"fcd00",-- -816
x"ffa00",-- -96
x"04300",-- 1072
x"05c00",-- 1472
x"05900",-- 1424
x"05800",-- 1408
x"06100",-- 1552
x"08f00",-- 2288
x"0cd00",-- 3280
x"0d700",-- 3440
x"0c600",-- 3168
x"0db00",-- 3504
x"0f100",-- 3856
x"13900",-- 5008
x"14400",-- 5184
x"0fd00",-- 4048
x"11200",-- 4384
x"15700",-- 5488
x"17000",-- 5888
x"18700",-- 6256
x"16700",-- 5744
x"14900",-- 5264
x"17a00",-- 6048
x"18d00",-- 6352
x"18500",-- 6224
x"14e00",-- 5344
x"11800",-- 4480
x"0fd00",-- 4048
x"0ee00",-- 3808
x"0c500",-- 3152
x"08100",-- 2064
x"04a00",-- 1184
x"fff00",-- -16
x"fb900",-- -1136
x"faf00",-- -1296
x"f8500",-- -1968
x"f4300",-- -3024
x"f2500",-- -3504
x"ef600",-- -4256
x"ed500",-- -4784
x"edf00",-- -4624
x"ee300",-- -4560
x"eae00",-- -5408
x"e8200",-- -6112
x"eab00",-- -5456
x"ecc00",-- -4928
x"ec300",-- -5072
x"eb700",-- -5264
x"ea800",-- -5504
x"ebb00",-- -5200
x"ef000",-- -4352
x"f0500",-- -4016
x"ee400",-- -4544
x"ee800",-- -4480
x"f1000",-- -3840
x"f2600",-- -3488
x"f4300",-- -3024
x"f4d00",-- -2864
x"f3900",-- -3184
x"f6200",-- -2528
x"f8500",-- -1968
x"f9700",-- -1680
x"fb300",-- -1232
x"fc500",-- -944
x"fd400",-- -704
x"fef00",-- -272
x"01a00",-- 416
x"02900",-- 656
x"03f00",-- 1008
x"05a00",-- 1440
x"05800",-- 1408
x"07900",-- 1936
x"09e00",-- 2528
x"0af00",-- 2800
x"0c100",-- 3088
x"0c800",-- 3200
x"0e600",-- 3680
x"10a00",-- 4256
x"14100",-- 5136
x"11600",-- 4448
x"0df00",-- 3568
x"13a00",-- 5024
x"17b00",-- 6064
x"16800",-- 5760
x"16600",-- 5728
x"14a00",-- 5280
x"15500",-- 5456
x"18f00",-- 6384
x"19100",-- 6416
x"16c00",-- 5824
x"12d00",-- 4816
x"11800",-- 4480
x"0ff00",-- 4080
x"0e200",-- 3616
x"0c800",-- 3200
x"07e00",-- 2016
x"02300",-- 560
x"feb00",-- -336
x"fd200",-- -736
x"fb400",-- -1216
x"f7900",-- -2160
x"f4500",-- -2992
x"f0f00",-- -3856
x"eed00",-- -4400
x"ef600",-- -4256
x"ef200",-- -4320
x"ed300",-- -4816
x"ead00",-- -5424
x"e9b00",-- -5712
x"e8b00",-- -5968
x"ebc00",-- -5184
x"f0800",-- -3968
x"ec500",-- -5040
x"e8e00",-- -5920
x"eb800",-- -5248
x"ed700",-- -4752
x"f1f00",-- -3600
x"f3800",-- -3200
x"ee300",-- -4560
x"ebd00",-- -5168
x"f1d00",-- -3632
x"f7600",-- -2208
x"f6500",-- -2480
x"f4e00",-- -2848
x"f4500",-- -2992
x"f5600",-- -2720
x"fb100",-- -1264
x"fe000",-- -512
x"fd400",-- -704
x"fc200",-- -992
x"fcf00",-- -784
x"01900",-- 400
x"05200",-- 1312
x"05800",-- 1408
x"04400",-- 1088
x"04800",-- 1152
x"06e00",-- 1760
x"09f00",-- 2544
x"0d700",-- 3440
x"0be00",-- 3040
x"0b000",-- 2816
x"0d900",-- 3472
x"11a00",-- 4512
x"14900",-- 5264
x"10400",-- 4160
x"0ee00",-- 3808
x"14200",-- 5152
x"15e00",-- 5600
x"16a00",-- 5792
x"16e00",-- 5856
x"14600",-- 5216
x"15f00",-- 5616
x"18000",-- 6144
x"17f00",-- 6128
x"15800",-- 5504
x"13200",-- 4896
x"10b00",-- 4272
x"0df00",-- 3568
x"0dc00",-- 3520
x"0a800",-- 2688
x"05c00",-- 1472
x"02600",-- 608
x"fd800",-- -640
x"fb800",-- -1152
x"fa700",-- -1424
x"f6900",-- -2416
x"f3300",-- -3280
x"f1500",-- -3760
x"efc00",-- -4160
x"ee200",-- -4576
x"eeb00",-- -4432
x"ee000",-- -4608
x"eb000",-- -5376
x"e9700",-- -5776
x"ea200",-- -5600
x"ee400",-- -4544
x"ef600",-- -4256
x"eb000",-- -5376
x"ea700",-- -5520
x"eca00",-- -4960
x"ef100",-- -4336
x"f3500",-- -3248
x"f1900",-- -3696
x"ec500",-- -5040
x"ef000",-- -4352
x"f5a00",-- -2656
x"f6a00",-- -2400
x"f5500",-- -2736
x"f5300",-- -2768
x"f4f00",-- -2832
x"f8500",-- -1968
x"fd300",-- -720
x"fd600",-- -672
x"fbf00",-- -1040
x"fcd00",-- -816
x"ffb00",-- -80
x"03900",-- 912
x"04d00",-- 1232
x"03e00",-- 992
x"04300",-- 1072
x"06700",-- 1648
x"08500",-- 2128
x"0ac00",-- 2752
x"0c800",-- 3200
x"0b400",-- 2880
x"0bc00",-- 3008
x"0f900",-- 3984
x"13f00",-- 5104
x"10300",-- 4144
x"0da00",-- 3488
x"13b00",-- 5040
x"16000",-- 5632
x"14300",-- 5168
x"15f00",-- 5616
x"15300",-- 5424
x"15800",-- 5504
x"18000",-- 6144
x"17300",-- 5936
x"15800",-- 5504
x"13800",-- 4992
x"12a00",-- 4768
x"0fe00",-- 4064
x"0d900",-- 3472
x"0b300",-- 2864
x"07700",-- 1904
x"04b00",-- 1200
x"00200",-- 32
x"fbd00",-- -1072
x"fae00",-- -1312
x"f8c00",-- -1856
x"f5400",-- -2752
x"f2000",-- -3584
x"f0700",-- -3984
x"ef800",-- -4224
x"ef100",-- -4336
x"eeb00",-- -4432
x"ebd00",-- -5168
x"e9f00",-- -5648
x"ebe00",-- -5152
x"ede00",-- -4640
x"ed200",-- -4832
x"ebc00",-- -5184
x"ebe00",-- -5152
x"edc00",-- -4672
x"ef200",-- -4320
x"f0400",-- -4032
x"f0600",-- -4000
x"eff00",-- -4112
x"f0700",-- -3984
x"f3100",-- -3312
x"f5200",-- -2784
x"f5100",-- -2800
x"f5500",-- -2736
x"f6300",-- -2512
x"f8400",-- -1984
x"fae00",-- -1312
x"fbe00",-- -1056
x"fc200",-- -992
x"fd700",-- -656
x"ffb00",-- -80
x"01500",-- 336
x"02700",-- 624
x"03600",-- 864
x"04400",-- 1088
x"05e00",-- 1504
x"07900",-- 1936
x"07d00",-- 2000
x"09400",-- 2368
x"0b100",-- 2832
x"0d100",-- 3344
x"0de00",-- 3552
x"0fb00",-- 4016
x"11300",-- 4400
x"0e500",-- 3664
x"10200",-- 4128
x"15200",-- 5408
x"15900",-- 5520
x"14600",-- 5216
x"14600",-- 5216
x"14900",-- 5264
x"16f00",-- 5872
x"17800",-- 6016
x"17100",-- 5904
x"14b00",-- 5296
x"11200",-- 4384
x"0fd00",-- 4048
x"0f800",-- 3968
x"0e400",-- 3648
x"09000",-- 2304
x"04d00",-- 1232
x"01b00",-- 432
x"fdc00",-- -576
x"fcc00",-- -832
x"fb600",-- -1184
x"f6900",-- -2416
x"f2300",-- -3536
x"f1600",-- -3744
x"f1700",-- -3728
x"f0600",-- -4000
x"ef300",-- -4304
x"ecd00",-- -4912
x"eb300",-- -5328
x"eba00",-- -5216
x"ed800",-- -4736
x"ee900",-- -4464
x"eca00",-- -4960
x"eb700",-- -5264
x"ed900",-- -4720
x"eeb00",-- -4432
x"f0000",-- -4096
x"f1600",-- -3744
x"f0b00",-- -3920
x"efe00",-- -4128
x"f1700",-- -3728
x"f4a00",-- -2912
x"f5c00",-- -2624
x"f6000",-- -2560
x"f6400",-- -2496
x"f6300",-- -2512
x"f8e00",-- -1824
x"fc500",-- -944
x"fdc00",-- -576
x"fd200",-- -736
x"fce00",-- -800
x"ff800",-- -128
x"02b00",-- 688
x"04700",-- 1136
x"04900",-- 1168
x"03d00",-- 976
x"04f00",-- 1264
x"07900",-- 1936
x"0b100",-- 2832
x"0bc00",-- 3008
x"0ac00",-- 2752
x"0ba00",-- 2976
x"0f000",-- 3840
x"12300",-- 4656
x"0f300",-- 3888
x"0eb00",-- 3760
x"13100",-- 4880
x"14f00",-- 5360
x"15100",-- 5392
x"14a00",-- 5280
x"13d00",-- 5072
x"16400",-- 5696
x"17f00",-- 6128
x"16d00",-- 5840
x"13d00",-- 5072
x"11f00",-- 4592
x"11500",-- 4432
x"0f900",-- 3984
x"0e300",-- 3632
x"09800",-- 2432
x"05500",-- 1360
x"03a00",-- 928
x"fff00",-- -16
x"fd100",-- -752
x"fab00",-- -1360
x"f7600",-- -2208
x"f4400",-- -3008
x"f2600",-- -3488
x"f2400",-- -3520
x"f0800",-- -3968
x"ee900",-- -4464
x"ed200",-- -4832
x"eca00",-- -4960
x"ecc00",-- -4928
x"ecf00",-- -4880
x"ede00",-- -4640
x"ecd00",-- -4912
x"eb800",-- -5248
x"ed900",-- -4720
x"ef500",-- -4272
x"ef800",-- -4224
x"ef900",-- -4208
x"efc00",-- -4160
x"f1400",-- -3776
x"f2200",-- -3552
x"f3700",-- -3216
x"f5500",-- -2736
x"f5200",-- -2784
x"f5900",-- -2672
x"f7e00",-- -2080
x"f9e00",-- -1568
x"fab00",-- -1360
x"fc200",-- -992
x"fd300",-- -720
x"fde00",-- -544
x"00800",-- 128
x"02d00",-- 720
x"02c00",-- 704
x"03700",-- 880
x"05000",-- 1280
x"06300",-- 1584
x"07900",-- 1936
x"09600",-- 2400
x"0ab00",-- 2736
x"0be00",-- 3040
x"0c500",-- 3152
x"0da00",-- 3488
x"10d00",-- 4304
x"0f300",-- 3888
x"0e000",-- 3584
x"12e00",-- 4832
x"15b00",-- 5552
x"13100",-- 4880
x"12500",-- 4688
x"14900",-- 5264
x"16f00",-- 5872
x"16300",-- 5680
x"15300",-- 5424
x"14000",-- 5120
x"11d00",-- 4560
x"10800",-- 4224
x"0f800",-- 3968
x"0e900",-- 3728
x"09d00",-- 2512
x"04b00",-- 1200
x"03a00",-- 928
x"00d00",-- 208
x"fd200",-- -736
x"fb300",-- -1232
x"f8100",-- -2032
x"f4400",-- -3008
x"f2c00",-- -3392
x"f2f00",-- -3344
x"f0900",-- -3952
x"eee00",-- -4384
x"eef00",-- -4368
x"ed200",-- -4832
x"ec500",-- -5040
x"ed500",-- -4784
x"ed800",-- -4736
x"edc00",-- -4672
x"ed800",-- -4736
x"ecf00",-- -4880
x"edf00",-- -4624
x"ef800",-- -4224
x"f0b00",-- -3920
x"f1a00",-- -3680
x"f1300",-- -3792
x"f0400",-- -4032
x"f3000",-- -3328
x"f6900",-- -2416
x"f6600",-- -2464
x"f6500",-- -2480
x"f7200",-- -2272
x"f8300",-- -2000
x"fb800",-- -1152
x"fe900",-- -368
x"fd500",-- -688
x"fcc00",-- -832
x"ffa00",-- -96
x"02500",-- 592
x"03a00",-- 928
x"04500",-- 1104
x"03f00",-- 1008
x"05400",-- 1344
x"07700",-- 1904
x"08f00",-- 2288
x"0ad00",-- 2768
x"0b900",-- 2960
x"0b200",-- 2848
x"0cf00",-- 3312
x"10d00",-- 4304
x"0ef00",-- 3824
x"0db00",-- 3504
x"12400",-- 4672
x"14700",-- 5232
x"13d00",-- 5072
x"13300",-- 4912
x"13100",-- 4880
x"15c00",-- 5568
x"17400",-- 5952
x"15e00",-- 5600
x"13600",-- 4960
x"11200",-- 4384
x"11200",-- 4384
x"10600",-- 4192
x"0e200",-- 3616
x"09e00",-- 2528
x"05a00",-- 1440
x"04400",-- 1088
x"01200",-- 288
x"fd500",-- -688
x"fba00",-- -1120
x"f9100",-- -1776
x"f5300",-- -2768
x"f2a00",-- -3424
x"f2300",-- -3536
x"f1400",-- -3776
x"f0800",-- -3968
x"eef00",-- -4368
x"ec000",-- -5120
x"ec700",-- -5008
x"edb00",-- -4688
x"ee000",-- -4608
x"ee700",-- -4496
x"ec700",-- -5008
x"eb800",-- -5248
x"eee00",-- -4384
x"f1100",-- -3824
x"f0700",-- -3984
x"ef200",-- -4320
x"f0900",-- -3952
x"f2700",-- -3472
x"f4100",-- -3056
x"f6300",-- -2512
x"f5c00",-- -2624
x"f5600",-- -2720
x"f8500",-- -1968
x"fb000",-- -1280
x"fbc00",-- -1088
x"fca00",-- -864
x"fd300",-- -720
x"fdd00",-- -560
x"00300",-- 48
x"03500",-- 848
x"03a00",-- 928
x"03800",-- 896
x"03d00",-- 976
x"04e00",-- 1248
x"07b00",-- 1968
x"0a300",-- 2608
x"09c00",-- 2496
x"09f00",-- 2544
x"0bd00",-- 3024
x"0dc00",-- 3520
x"10300",-- 4144
x"0e900",-- 3728
x"0d900",-- 3472
x"11500",-- 4432
x"14f00",-- 5360
x"14400",-- 5184
x"11b00",-- 4528
x"11e00",-- 4576
x"17100",-- 5904
x"17900",-- 6032
x"14800",-- 5248
x"12a00",-- 4768
x"11300",-- 4400
x"11600",-- 4448
x"10700",-- 4208
x"0d700",-- 3440
x"08a00",-- 2208
x"05f00",-- 1520
x"04400",-- 1088
x"01100",-- 272
x"fda00",-- -608
x"fac00",-- -1344
x"f8800",-- -1920
x"f6000",-- -2560
x"f2f00",-- -3344
x"f1d00",-- -3632
x"f1d00",-- -3632
x"f0200",-- -4064
x"ee100",-- -4592
x"ed100",-- -4848
x"ed100",-- -4848
x"edb00",-- -4688
x"eec00",-- -4416
x"eda00",-- -4704
x"ebb00",-- -5200
x"ed200",-- -4832
x"efb00",-- -4176
x"f0000",-- -4096
x"ef900",-- -4208
x"f0400",-- -4032
x"f1200",-- -3808
x"f2b00",-- -3408
x"f5200",-- -2784
x"f5e00",-- -2592
x"f5c00",-- -2624
x"f6d00",-- -2352
x"f9200",-- -1760
x"fb300",-- -1232
x"fcb00",-- -848
x"fcd00",-- -816
x"fd000",-- -768
x"ff900",-- -112
x"02000",-- 512
x"02400",-- 576
x"02600",-- 608
x"04000",-- 1024
x"05600",-- 1376
x"06100",-- 1552
x"07c00",-- 1984
x"09400",-- 2368
x"09700",-- 2416
x"0bb00",-- 2992
x"0cb00",-- 3248
x"0d700",-- 3440
x"0ed00",-- 3792
x"0de00",-- 3552
x"0ed00",-- 3792
x"12000",-- 4608
x"13700",-- 4976
x"14700",-- 5232
x"12900",-- 4752
x"10c00",-- 4288
x"14f00",-- 5360
x"18300",-- 6192
x"16300",-- 5680
x"10200",-- 4128
x"0e900",-- 3728
x"0fb00",-- 4016
x"0ff00",-- 4080
x"0fb00",-- 4016
x"09600",-- 2400
x"01900",-- 400
x"fff00",-- -16
x"00b00",-- 176
x"00000",-- 0
x"fbc00",-- -1088
x"f5d00",-- -2608
x"f2400",-- -3520
x"f1900",-- -3696
x"f4100",-- -3056
x"f3700",-- -3216
x"ef500",-- -4272
x"eb900",-- -5232
x"eb700",-- -5264
x"ee000",-- -4608
x"eff00",-- -4112
x"ef800",-- -4224
x"ec700",-- -5008
x"eb300",-- -5328
x"edf00",-- -4624
x"f0f00",-- -3856
x"f1a00",-- -3680
x"f0200",-- -4064
x"eff00",-- -4112
x"f1a00",-- -3680
x"f3f00",-- -3088
x"f7500",-- -2224
x"f7d00",-- -2096
x"f6600",-- -2464
x"f6e00",-- -2336
x"f9c00",-- -1600
x"fd800",-- -640
x"fdf00",-- -528
x"fd400",-- -704
x"fdb00",-- -592
x"ff100",-- -240
x"01e00",-- 480
x"04100",-- 1040
x"04600",-- 1120
x"03700",-- 880
x"03f00",-- 1008
x"06a00",-- 1696
x"08a00",-- 2208
x"09400",-- 2368
x"0a600",-- 2656
x"0b500",-- 2896
x"0b500",-- 2896
x"0d800",-- 3456
x"0ea00",-- 3744
x"0df00",-- 3568
x"10d00",-- 4304
x"12500",-- 4688
x"10700",-- 4208
x"11500",-- 4432
x"13b00",-- 5040
x"15400",-- 5440
x"15600",-- 5472
x"13a00",-- 5024
x"13700",-- 4976
x"11700",-- 4464
x"10b00",-- 4272
x"10200",-- 4128
x"0d900",-- 3472
x"0a800",-- 2688
x"06f00",-- 1776
x"03f00",-- 1008
x"02c00",-- 704
x"00800",-- 128
x"fc300",-- -976
x"f8600",-- -1952
x"f7500",-- -2224
x"f4f00",-- -2832
x"f3800",-- -3200
x"f4800",-- -2944
x"efe00",-- -4128
x"ecf00",-- -4880
x"efb00",-- -4176
x"f0600",-- -4000
x"ee900",-- -4464
x"ed700",-- -4752
x"ec200",-- -5088
x"ec700",-- -5008
x"ef900",-- -4208
x"f0b00",-- -3920
x"ee500",-- -4528
x"edf00",-- -4624
x"efe00",-- -4128
x"f2b00",-- -3408
x"f4c00",-- -2880
x"f4900",-- -2928
x"f4000",-- -3072
x"f4a00",-- -2912
x"f7a00",-- -2144
x"faf00",-- -1296
x"fb400",-- -1216
x"fa800",-- -1408
x"fa700",-- -1424
x"fd100",-- -752
x"00700",-- 112
x"01a00",-- 416
x"01100",-- 272
x"00c00",-- 192
x"02c00",-- 704
x"05400",-- 1344
x"06700",-- 1648
x"06d00",-- 1744
x"07a00",-- 1952
x"09500",-- 2384
x"0af00",-- 2800
x"0c000",-- 3072
x"0cf00",-- 3312
x"0ef00",-- 3824
x"0de00",-- 3552
x"0cb00",-- 3248
x"0f600",-- 3936
x"12f00",-- 4848
x"14500",-- 5200
x"12f00",-- 4848
x"11800",-- 4480
x"13700",-- 4976
x"14e00",-- 5344
x"14100",-- 5136
x"13400",-- 4928
x"12100",-- 4624
x"10900",-- 4240
x"0d200",-- 3360
x"0a600",-- 2656
x"09700",-- 2416
x"08d00",-- 2256
x"05b00",-- 1456
x"00000",-- 0
x"fb800",-- -1152
x"f9f00",-- -1552
x"fab00",-- -1360
x"f9d00",-- -1584
x"f4800",-- -2944
x"f1300",-- -3792
x"f0000",-- -4096
x"f0700",-- -3984
x"f1200",-- -3808
x"efa00",-- -4192
x"ed200",-- -4832
x"ece00",-- -4896
x"ed400",-- -4800
x"ed700",-- -4752
x"eea00",-- -4448
x"eee00",-- -4384
x"ee100",-- -4592
x"ed300",-- -4816
x"ef300",-- -4304
x"f2300",-- -3536
x"f2f00",-- -3344
x"f3800",-- -3200
x"f4200",-- -3040
x"f3e00",-- -3104
x"f7600",-- -2208
x"fb100",-- -1264
x"fa600",-- -1440
x"f9f00",-- -1552
x"fbb00",-- -1104
x"fcc00",-- -832
x"ff200",-- -224
x"02a00",-- 672
x"01900",-- 400
x"ffb00",-- -80
x"02700",-- 624
x"05500",-- 1360
x"06700",-- 1648
x"06b00",-- 1712
x"06000",-- 1536
x"06f00",-- 1776
x"0a100",-- 2576
x"0c900",-- 3216
x"0c100",-- 3088
x"0bd00",-- 3024
x"0ea00",-- 3744
x"0dc00",-- 3520
x"0e200",-- 3616
x"11500",-- 4432
x"12f00",-- 4848
x"13200",-- 4896
x"12300",-- 4656
x"11700",-- 4464
x"13800",-- 4992
x"15a00",-- 5536
x"15600",-- 5472
x"12a00",-- 4768
x"0f100",-- 3856
x"0d600",-- 3424
x"0d700",-- 3440
x"0de00",-- 3552
x"0a100",-- 2576
x"03c00",-- 960
x"ffd00",-- -48
x"ff300",-- -208
x"fe900",-- -368
x"fc000",-- -1024
x"f7a00",-- -2144
x"f2a00",-- -3424
x"f2000",-- -3584
x"f3200",-- -3296
x"f1b00",-- -3664
x"ef500",-- -4272
x"ecd00",-- -4912
x"ec400",-- -5056
x"edb00",-- -4688
x"ee900",-- -4464
x"ed200",-- -4832
x"eba00",-- -5216
x"ecf00",-- -4880
x"ed800",-- -4736
x"ee400",-- -4544
x"f0600",-- -4000
x"efb00",-- -4176
x"f0900",-- -3952
x"f3800",-- -3200
x"f4500",-- -2992
x"f4d00",-- -2864
x"f7700",-- -2192
x"f9200",-- -1760
x"f9a00",-- -1632
x"fb400",-- -1216
x"fc700",-- -912
x"fcb00",-- -848
x"ff600",-- -160
x"01400",-- 320
x"00900",-- 144
x"00d00",-- 208
x"02e00",-- 736
x"05700",-- 1392
x"05c00",-- 1472
x"05d00",-- 1488
x"06200",-- 1568
x"08100",-- 2064
x"0ad00",-- 2768
x"0af00",-- 2800
x"0b700",-- 2928
x"0be00",-- 3040
x"0e500",-- 3664
x"0df00",-- 3568
x"0d900",-- 3472
x"10800",-- 4224
x"12100",-- 4624
x"12b00",-- 4784
x"12e00",-- 4832
x"11b00",-- 4528
x"12200",-- 4640
x"14800",-- 5248
x"16000",-- 5632
x"14600",-- 5216
x"0ed00",-- 3792
x"0cf00",-- 3312
x"0d900",-- 3472
x"0e700",-- 3696
x"0c200",-- 3104
x"05300",-- 1328
x"ff800",-- -128
x"fee00",-- -288
x"ffb00",-- -80
x"fde00",-- -544
x"f8200",-- -2016
x"f3100",-- -3312
x"f2100",-- -3568
x"f2700",-- -3472
x"f2700",-- -3472
x"f0b00",-- -3920
x"ecd00",-- -4912
x"eb700",-- -5264
x"ed000",-- -4864
x"ee300",-- -4560
x"ed800",-- -4736
x"ec000",-- -5120
x"ebd00",-- -5168
x"ecf00",-- -4880
x"ee800",-- -4480
x"ef700",-- -4240
x"eff00",-- -4112
x"f0100",-- -4080
x"f2500",-- -3504
x"f4e00",-- -2848
x"f5800",-- -2688
x"f6000",-- -2560
x"f7b00",-- -2128
x"f9e00",-- -1568
x"fc100",-- -1008
x"fcd00",-- -816
x"fc300",-- -976
x"fdb00",-- -592
x"00f00",-- 240
x"02100",-- 528
x"01f00",-- 496
x"02600",-- 608
x"03400",-- 832
x"05400",-- 1344
x"06f00",-- 1776
x"07900",-- 1936
x"07b00",-- 1968
x"08300",-- 2096
x"0a800",-- 2688
x"0d500",-- 3408
x"0c500",-- 3152
x"0ce00",-- 3296
x"0ec00",-- 3776
x"0dd00",-- 3536
x"0ff00",-- 4080
x"12400",-- 4672
x"12b00",-- 4784
x"12a00",-- 4768
x"13d00",-- 5072
x"13600",-- 4960
x"13600",-- 4960
x"14800",-- 5248
x"15c00",-- 5568
x"12900",-- 4752
x"0e100",-- 3600
x"0ca00",-- 3232
x"0d200",-- 3360
x"0c400",-- 3136
x"08100",-- 2064
x"02d00",-- 720
x"fe800",-- -384
x"fd100",-- -752
x"fc600",-- -928
x"fa100",-- -1520
x"f6100",-- -2544
x"f2300",-- -3536
x"f0300",-- -4048
x"eff00",-- -4112
x"efe00",-- -4128
x"ef100",-- -4336
x"ecc00",-- -4928
x"eb700",-- -5264
x"eb500",-- -5296
x"ebf00",-- -5136
x"eca00",-- -4960
x"ed200",-- -4832
x"ecf00",-- -4880
x"ec800",-- -4992
x"ed800",-- -4736
x"efd00",-- -4144
x"f1900",-- -3696
x"f3000",-- -3328
x"f3900",-- -3184
x"f4300",-- -3024
x"f6400",-- -2496
x"f8900",-- -1904
x"fa700",-- -1424
x"fc200",-- -992
x"fcb00",-- -848
x"fc900",-- -880
x"fe700",-- -400
x"01500",-- 336
x"02800",-- 640
x"02500",-- 592
x"02b00",-- 688
x"03d00",-- 976
x"05a00",-- 1440
x"07700",-- 1904
x"07d00",-- 2000
x"07f00",-- 2032
x"09a00",-- 2464
x"0b700",-- 2928
x"0cc00",-- 3264
x"0cc00",-- 3264
x"0dc00",-- 3520
x"10c00",-- 4288
x"0e800",-- 3712
x"0e900",-- 3728
x"12300",-- 4656
x"14800",-- 5248
x"15300",-- 5424
x"13e00",-- 5088
x"11d00",-- 4560
x"12e00",-- 4832
x"16500",-- 5712
x"16f00",-- 5872
x"13300",-- 4912
x"0e900",-- 3728
x"0bc00",-- 3008
x"0c000",-- 3072
x"0cd00",-- 3280
x"09600",-- 2400
x"03000",-- 768
x"fd900",-- -624
x"fb500",-- -1200
x"fb100",-- -1264
x"fa700",-- -1424
x"f6e00",-- -2336
x"f1300",-- -3792
x"edf00",-- -4624
x"ee600",-- -4512
x"ee700",-- -4496
x"ef500",-- -4272
x"ecf00",-- -4880
x"e9700",-- -5776
x"e8e00",-- -5920
x"eb600",-- -5280
x"ecd00",-- -4912
x"ec600",-- -5024
x"ec400",-- -5056
x"eaf00",-- -5392
x"ed200",-- -4832
x"f0c00",-- -3904
x"f1500",-- -3760
x"f1d00",-- -3632
x"f4100",-- -3056
x"f4e00",-- -2848
x"f6800",-- -2432
x"f9300",-- -1744
x"fa800",-- -1408
x"fba00",-- -1120
x"fd900",-- -624
x"fe400",-- -448
x"ff100",-- -240
x"01b00",-- 432
x"02f00",-- 752
x"03400",-- 832
x"04300",-- 1072
x"04d00",-- 1232
x"06200",-- 1568
x"07a00",-- 1952
x"09600",-- 2400
x"09e00",-- 2528
x"0ab00",-- 2736
x"0b900",-- 2960
x"0ce00",-- 3296
x"0e900",-- 3728
x"0ff00",-- 4080
x"0fd00",-- 4048
x"0e600",-- 3680
x"10700",-- 4208
x"12e00",-- 4832
x"15100",-- 5392
x"15500",-- 5456
x"13700",-- 4976
x"12700",-- 4720
x"13f00",-- 5104
x"15e00",-- 5600
x"15b00",-- 5552
x"12400",-- 4672
x"0e100",-- 3600
x"0b600",-- 2912
x"0b800",-- 2944
x"0b700",-- 2928
x"07f00",-- 2032
x"01600",-- 352
x"fc400",-- -960
x"fa100",-- -1520
x"f9f00",-- -1552
x"f9c00",-- -1600
x"f4c00",-- -2880
x"eea00",-- -4448
x"ec400",-- -5056
x"ed700",-- -4752
x"ef300",-- -4304
x"ee200",-- -4576
x"ea900",-- -5488
x"e7d00",-- -6192
x"e7f00",-- -6160
x"eb200",-- -5344
x"ed300",-- -4816
x"ed300",-- -4816
x"ea800",-- -5504
x"e9d00",-- -5680
x"eda00",-- -4704
x"f1500",-- -3760
x"f3c00",-- -3136
x"f3f00",-- -3088
x"f2b00",-- -3408
x"f3c00",-- -3136
x"f7500",-- -2224
x"fb500",-- -1200
x"fd600",-- -672
x"fcd00",-- -816
x"fc000",-- -1024
x"fd700",-- -656
x"01900",-- 400
x"04200",-- 1056
x"03b00",-- 944
x"03900",-- 912
x"04e00",-- 1248
x"05e00",-- 1504
x"06d00",-- 1744
x"08500",-- 2128
x"09600",-- 2400
x"0ad00",-- 2768
x"0b400",-- 2880
x"0b200",-- 2848
x"0d200",-- 3360
x"0ea00",-- 3744
x"11c00",-- 4544
x"11100",-- 4368
x"0e000",-- 3584
x"10000",-- 4096
x"13f00",-- 5104
x"16a00",-- 5792
x"16300",-- 5680
x"13400",-- 4928
x"11d00",-- 4560
x"14100",-- 5136
x"16b00",-- 5808
x"16700",-- 5744
x"12000",-- 4608
x"0c400",-- 3136
x"09b00",-- 2480
x"0b500",-- 2896
x"0af00",-- 2800
x"06500",-- 1616
x"ff300",-- -208
x"f9900",-- -1648
x"f8200",-- -2016
x"f9000",-- -1792
x"f7700",-- -2192
x"f1900",-- -3696
x"ec700",-- -5008
x"eae00",-- -5408
x"ec400",-- -5056
x"ee300",-- -4560
x"ebe00",-- -5152
x"e8200",-- -6112
x"e6d00",-- -6448
x"e9100",-- -5872
x"eb800",-- -5248
x"ebd00",-- -5168
x"ea800",-- -5504
x"ea000",-- -5632
x"ec600",-- -5024
x"ef900",-- -4208
x"f2100",-- -3568
x"f2900",-- -3440
x"f2500",-- -3504
x"f3800",-- -3200
x"f7500",-- -2224
x"fa500",-- -1456
x"fb100",-- -1264
x"fb800",-- -1152
x"fc400",-- -960
x"fea00",-- -352
x"02500",-- 592
x"03600",-- 864
x"03100",-- 784
x"03800",-- 896
x"05500",-- 1360
x"07700",-- 1904
x"09000",-- 2304
x"08300",-- 2096
x"08700",-- 2160
x"0aa00",-- 2720
x"0ce00",-- 3296
x"0d700",-- 3440
x"0e700",-- 3696
x"0e200",-- 3616
x"10300",-- 4144
x"13100",-- 4880
x"10900",-- 4240
x"10300",-- 4144
x"11b00",-- 4528
x"15a00",-- 5536
x"17400",-- 5952
x"15f00",-- 5616
x"12100",-- 4624
x"11a00",-- 4512
x"14400",-- 5184
x"17400",-- 5952
x"15000",-- 5376
x"0e400",-- 3648
x"08d00",-- 2256
x"07c00",-- 1984
x"09f00",-- 2544
x"08e00",-- 2272
x"03500",-- 848
x"fa800",-- -1408
x"f5900",-- -2672
x"f5c00",-- -2624
x"f7100",-- -2288
x"f4e00",-- -2848
x"ef200",-- -4320
x"e9400",-- -5824
x"e8200",-- -6112
x"eb500",-- -5296
x"eca00",-- -4960
x"ea800",-- -5504
x"e7600",-- -6304
x"e6500",-- -6576
x"e8300",-- -6096
x"eb200",-- -5344
x"eb700",-- -5264
x"eb000",-- -5376
x"ec600",-- -5024
x"ee000",-- -4608
x"f0700",-- -3984
x"f1f00",-- -3600
x"f2c00",-- -3392
x"f5000",-- -2816
x"f7b00",-- -2128
x"f9000",-- -1792
x"f9f00",-- -1552
x"fb500",-- -1200
x"fd400",-- -704
x"00100",-- 16
x"02c00",-- 704
x"03300",-- 816
x"03400",-- 832
x"04900",-- 1168
x"06a00",-- 1696
x"09500",-- 2384
x"0ac00",-- 2752
x"09700",-- 2416
x"09200",-- 2336
x"0b600",-- 2912
x"0e600",-- 3680
x"0f900",-- 3984
x"10300",-- 4144
x"0fb00",-- 4016
x"10a00",-- 4256
x"14400",-- 5184
x"11e00",-- 4576
x"11800",-- 4480
x"12e00",-- 4832
x"15400",-- 5440
x"17300",-- 5936
x"15f00",-- 5616
x"12900",-- 4752
x"11200",-- 4384
x"13b00",-- 5040
x"15f00",-- 5616
x"13f00",-- 5104
x"0e800",-- 3712
x"08100",-- 2064
x"05c00",-- 1472
x"08100",-- 2064
x"07700",-- 1904
x"02900",-- 656
x"fa300",-- -1488
x"f4000",-- -3072
x"f3200",-- -3296
x"f4800",-- -2944
x"f3800",-- -3200
x"ede00",-- -4640
x"e8300",-- -6096
x"e7600",-- -6304
x"e8800",-- -6016
x"eaa00",-- -5472
x"e9b00",-- -5712
x"e7300",-- -6352
x"e6200",-- -6624
x"e8000",-- -6144
x"e9e00",-- -5664
x"ea100",-- -5616
x"ebb00",-- -5200
x"ed000",-- -4864
x"ee900",-- -4464
x"f1900",-- -3696
x"f2a00",-- -3424
x"f2e00",-- -3360
x"f5c00",-- -2624
x"f8c00",-- -1856
x"fb000",-- -1280
x"fc400",-- -960
x"fc600",-- -928
x"fce00",-- -800
x"fff00",-- -16
x"04100",-- 1040
x"05400",-- 1344
x"04900",-- 1168
x"04b00",-- 1200
x"06c00",-- 1728
x"09d00",-- 2512
x"0b900",-- 2960
x"0a900",-- 2704
x"09500",-- 2384
x"0b900",-- 2960
x"0ed00",-- 3792
x"0f900",-- 3984
x"0fd00",-- 4048
x"0f700",-- 3952
x"11200",-- 4384
x"13900",-- 5008
x"11700",-- 4464
x"10f00",-- 4336
x"11a00",-- 4512
x"14b00",-- 5296
x"17600",-- 5984
x"15d00",-- 5584
x"12200",-- 4640
x"10600",-- 4192
x"11d00",-- 4560
x"15200",-- 5408
x"14a00",-- 5280
x"0ef00",-- 3824
x"07d00",-- 2000
x"04800",-- 1152
x"06100",-- 1552
x"06700",-- 1648
x"03200",-- 800
x"fb100",-- -1264
x"f3a00",-- -3168
x"f1b00",-- -3664
x"f2800",-- -3456
x"f2c00",-- -3392
x"ee900",-- -4464
x"e9d00",-- -5680
x"e7000",-- -6400
x"e7100",-- -6384
x"e8900",-- -6000
x"e8300",-- -6096
x"e7e00",-- -6176
x"e7100",-- -6384
x"e7e00",-- -6176
x"e8900",-- -6000
x"e8700",-- -6032
x"ea700",-- -5520
x"ed300",-- -4816
x"f0000",-- -4096
x"f1c00",-- -3648
x"f1900",-- -3696
x"f1a00",-- -3680
x"f4b00",-- -2896
x"f9400",-- -1728
x"fbf00",-- -1040
x"fc100",-- -1008
x"fbf00",-- -1040
x"fce00",-- -800
x"ffd00",-- -48
x"04500",-- 1104
x"06800",-- 1664
x"05b00",-- 1456
x"05300",-- 1328
x"07700",-- 1904
x"0a700",-- 2672
x"0ca00",-- 3232
x"0c600",-- 3168
x"0c400",-- 3136
x"0d100",-- 3344
x"0f800",-- 3968
x"11b00",-- 4528
x"12500",-- 4688
x"12200",-- 4640
x"15400",-- 5440
x"15600",-- 5472
x"12c00",-- 4800
x"13400",-- 4928
x"14000",-- 5120
x"17c00",-- 6080
x"19800",-- 6528
x"16b00",-- 5808
x"12100",-- 4624
x"10c00",-- 4288
x"12d00",-- 4816
x"14f00",-- 5360
x"12d00",-- 4816
x"0d200",-- 3360
x"05900",-- 1424
x"02800",-- 640
x"03e00",-- 992
x"03100",-- 784
x"fec00",-- -320
x"f7900",-- -2160
x"f1900",-- -3696
x"ee600",-- -4512
x"ef000",-- -4352
x"edd00",-- -4656
x"eb000",-- -5376
x"e7d00",-- -6192
x"e6400",-- -6592
x"e5400",-- -6848
x"e5000",-- -6912
x"e5900",-- -6768
x"e6100",-- -6640
x"e7d00",-- -6192
x"e8f00",-- -5904
x"e8b00",-- -5968
x"e7c00",-- -6208
x"ea300",-- -5584
x"ee200",-- -4576
x"f2200",-- -3552
x"f4300",-- -3024
x"f3800",-- -3200
x"f3200",-- -3296
x"f5e00",-- -2592
x"fa800",-- -1408
x"fe200",-- -480
x"ff000",-- -256
x"ff000",-- -256
x"ff400",-- -192
x"01200",-- 288
x"04f00",-- 1264
x"07700",-- 1904
x"07d00",-- 2000
x"08500",-- 2128
x"09500",-- 2384
x"0a800",-- 2688
x"0bd00",-- 3024
x"0cd00",-- 3280
x"0e100",-- 3600
x"10800",-- 4224
x"11200",-- 4384
x"11c00",-- 4544
x"11400",-- 4416
x"14400",-- 5184
x"16e00",-- 5856
x"13a00",-- 5024
x"14000",-- 5120
x"13600",-- 4960
x"16600",-- 5728
x"18000",-- 6144
x"17d00",-- 6096
x"12500",-- 4688
x"0ea00",-- 3744
x"11800",-- 4480
x"13a00",-- 5024
x"15000",-- 5376
x"0f500",-- 3920
x"05900",-- 1424
x"00600",-- 96
x"01700",-- 368
x"03800",-- 896
x"00600",-- 96
x"f9400",-- -1728
x"f0c00",-- -3904
x"ebb00",-- -5200
x"ee100",-- -4592
x"eed00",-- -4400
x"eca00",-- -4960
x"e9600",-- -5792
x"e6000",-- -6656
x"e5000",-- -6912
x"e6200",-- -6624
x"e6e00",-- -6432
x"e7800",-- -6272
x"e9700",-- -5776
x"ec100",-- -5104
x"eb000",-- -5376
x"ea300",-- -5584
x"ea800",-- -5504
x"ed700",-- -4752
x"f3900",-- -3184
x"f7c00",-- -2112
x"f7100",-- -2288
x"f4500",-- -2992
x"f5400",-- -2752
x"f9000",-- -1792
x"feb00",-- -336
x"02600",-- 608
x"01000",-- 256
x"fe700",-- -400
x"ffd00",-- -48
x"03700",-- 880
x"06c00",-- 1728
x"08500",-- 2128
x"08000",-- 2048
x"07b00",-- 1968
x"08900",-- 2192
x"0a400",-- 2624
x"0a700",-- 2672
x"0ba00",-- 2976
x"0df00",-- 3568
x"0ee00",-- 3808
x"0f800",-- 3968
x"10300",-- 4144
x"10500",-- 4176
x"13900",-- 5008
x"13600",-- 4960
x"13200",-- 4896
x"12e00",-- 4832
x"13200",-- 4896
x"16200",-- 5664
x"16400",-- 5696
x"15500",-- 5456
x"13300",-- 4912
x"12300",-- 4656
x"12200",-- 4640
x"12700",-- 4720
x"10700",-- 4208
x"0c600",-- 3168
x"06d00",-- 1744
x"04700",-- 1136
x"03200",-- 800
x"01000",-- 256
x"fda00",-- -608
x"f7900",-- -2160
x"f3300",-- -3280
x"f0c00",-- -3904
x"ef600",-- -4256
x"ee500",-- -4528
x"eb200",-- -5344
x"e9b00",-- -5712
x"e7b00",-- -6224
x"e7900",-- -6256
x"e7c00",-- -6208
x"e6d00",-- -6448
x"e7c00",-- -6208
x"e8900",-- -6000
x"ea900",-- -5488
x"ea800",-- -5504
x"eb000",-- -5376
x"ebf00",-- -5136
x"ee700",-- -4496
x"f2400",-- -3520
x"f4b00",-- -2896
x"f4b00",-- -2896
x"f5500",-- -2736
x"f6e00",-- -2336
x"f9800",-- -1664
x"fd000",-- -768
x"ff100",-- -240
x"ffa00",-- -96
x"fff00",-- -16
x"02200",-- 544
x"04200",-- 1056
x"05a00",-- 1440
x"06d00",-- 1744
x"07a00",-- 1952
x"08f00",-- 2288
x"0a200",-- 2592
x"0b000",-- 2816
x"0b100",-- 2832
x"0ba00",-- 2976
x"0d800",-- 3456
x"0e500",-- 3664
x"10400",-- 4160
x"10a00",-- 4256
x"11500",-- 4432
x"13d00",-- 5072
x"11b00",-- 4528
x"12000",-- 4608
x"12a00",-- 4768
x"14000",-- 5120
x"16800",-- 5760
x"16000",-- 5632
x"13600",-- 4960
x"11d00",-- 4560
x"10c00",-- 4288
x"11d00",-- 4560
x"12300",-- 4656
x"0f800",-- 3968
x"0b900",-- 2960
x"05b00",-- 1456
x"03d00",-- 976
x"02100",-- 528
x"fff00",-- -16
x"fd600",-- -672
x"f8000",-- -2048
x"f3e00",-- -3104
x"f0e00",-- -3872
x"ee900",-- -4464
x"ed100",-- -4848
x"ebd00",-- -5168
x"eae00",-- -5408
x"e9800",-- -5760
x"e8900",-- -6000
x"e7100",-- -6384
x"e6300",-- -6608
x"e8000",-- -6144
x"e9e00",-- -5664
x"eb200",-- -5344
x"eba00",-- -5216
x"eb400",-- -5312
x"ec100",-- -5104
x"ee800",-- -4480
x"f2500",-- -3504
x"f4400",-- -3008
x"f5300",-- -2768
x"f6d00",-- -2352
x"f8000",-- -2048
x"fa500",-- -1456
x"fcb00",-- -848
x"fd900",-- -624
x"ff400",-- -192
x"01800",-- 384
x"03e00",-- 992
x"04000",-- 1024
x"04b00",-- 1200
x"05d00",-- 1488
x"07400",-- 1856
x"08b00",-- 2224
x"0aa00",-- 2720
x"0a800",-- 2688
x"09500",-- 2384
x"0a700",-- 2672
x"0b500",-- 2896
x"0e900",-- 3728
x"0eb00",-- 3760
x"0f700",-- 3952
x"10300",-- 4144
x"12200",-- 4640
x"11100",-- 4368
x"10000",-- 4096
x"11700",-- 4464
x"11d00",-- 4560
x"15d00",-- 5584
x"16300",-- 5680
x"13e00",-- 5088
x"10e00",-- 4320
x"0f800",-- 3968
x"10e00",-- 4320
x"11700",-- 4464
x"10d00",-- 4304
x"0d600",-- 3424
x"07600",-- 1888
x"04900",-- 1168
x"03000",-- 768
x"00e00",-- 224
x"feb00",-- -336
x"fa600",-- -1440
x"f6c00",-- -2368
x"f3b00",-- -3152
x"f1600",-- -3744
x"ef600",-- -4256
x"eca00",-- -4960
x"ec500",-- -5040
x"eba00",-- -5216
x"eb200",-- -5344
x"ea500",-- -5552
x"e8200",-- -6112
x"e8000",-- -6144
x"e9000",-- -5888
x"ebb00",-- -5200
x"ec500",-- -5040
x"ece00",-- -4896
x"ed700",-- -4752
x"ee600",-- -4512
x"f0e00",-- -3872
x"f3600",-- -3232
x"f4b00",-- -2896
x"f6400",-- -2496
x"f8500",-- -1968
x"f9e00",-- -1568
x"fb900",-- -1136
x"fd100",-- -752
x"fe900",-- -368
x"ff900",-- -112
x"02000",-- 512
x"03a00",-- 928
x"04400",-- 1088
x"04700",-- 1136
x"05d00",-- 1488
x"06300",-- 1584
x"08900",-- 2192
x"09900",-- 2448
x"07e00",-- 2016
x"09000",-- 2304
x"09a00",-- 2464
x"0b800",-- 2944
x"0bc00",-- 3008
x"0c400",-- 3136
x"0d400",-- 3392
x"0e500",-- 3664
x"11800",-- 4480
x"10e00",-- 4320
x"0fb00",-- 4016
x"0f400",-- 3904
x"10b00",-- 4272
x"13000",-- 4864
x"14500",-- 5200
x"13600",-- 4960
x"10b00",-- 4272
x"10500",-- 4176
x"0fd00",-- 4048
x"0ff00",-- 4080
x"0e900",-- 3728
x"0c500",-- 3152
x"08c00",-- 2240
x"06800",-- 1664
x"04e00",-- 1248
x"01700",-- 368
x"feb00",-- -336
x"fa700",-- -1424
x"f8e00",-- -1824
x"f6700",-- -2448
x"f4a00",-- -2912
x"f1b00",-- -3664
x"ee200",-- -4576
x"ed900",-- -4720
x"ecf00",-- -4880
x"ed300",-- -4816
x"ec300",-- -5072
x"eac00",-- -5440
x"e9d00",-- -5680
x"eb000",-- -5376
x"ec100",-- -5104
x"ed000",-- -4864
x"ed900",-- -4720
x"ee000",-- -4608
x"efb00",-- -4176
x"f1a00",-- -3680
x"f3b00",-- -3152
x"f4500",-- -2992
x"f5c00",-- -2624
x"f7c00",-- -2112
x"f9e00",-- -1568
x"fb800",-- -1152
x"fc800",-- -896
x"fdb00",-- -592
x"fed00",-- -304
x"00a00",-- 160
x"02200",-- 544
x"02400",-- 576
x"03d00",-- 976
x"04b00",-- 1200
x"03c00",-- 960
x"07600",-- 1888
x"06100",-- 1552
x"05600",-- 1376
x"06600",-- 1632
x"08700",-- 2160
x"08d00",-- 2256
x"08e00",-- 2272
x"0c100",-- 3088
x"09100",-- 2320
x"0cb00",-- 3248
x"0ce00",-- 3296
x"0f200",-- 3872
x"0f800",-- 3968
x"0e700",-- 3696
x"0f900",-- 3984
x"0f100",-- 3856
x"12500",-- 4688
x"12700",-- 4720
x"11d00",-- 4560
x"0fa00",-- 4000
x"10900",-- 4240
x"0f000",-- 3840
x"0f600",-- 3936
x"0db00",-- 3504
x"0b700",-- 2928
x"09200",-- 2336
x"06b00",-- 1712
x"05e00",-- 1504
x"01800",-- 384
x"ffb00",-- -80
x"fc300",-- -976
x"fa400",-- -1472
x"f8100",-- -2032
x"f6700",-- -2448
x"f3700",-- -3216
x"f1200",-- -3808
x"f0a00",-- -3936
x"efb00",-- -4176
x"ef800",-- -4224
x"edc00",-- -4672
x"ed800",-- -4736
x"ec200",-- -5088
x"edd00",-- -4656
x"ee300",-- -4560
x"ee200",-- -4576
x"eea00",-- -4448
x"eef00",-- -4368
x"f1500",-- -3760
x"f2800",-- -3456
x"f4800",-- -2944
x"f5000",-- -2816
x"f5800",-- -2688
x"f7600",-- -2208
x"f9000",-- -1792
x"fac00",-- -1344
x"fc300",-- -976
x"fd300",-- -720
x"fd600",-- -672
x"fe600",-- -416
x"01900",-- 400
x"ffb00",-- -80
x"01700",-- 368
x"03400",-- 832
x"02700",-- 624
x"04300",-- 1072
x"04300",-- 1072
x"03f00",-- 1008
x"02800",-- 640
x"06f00",-- 1776
x"06c00",-- 1728
x"05700",-- 1392
x"08200",-- 2080
x"07700",-- 1904
x"09100",-- 2320
x"0b000",-- 2816
x"0a800",-- 2688
x"0c800",-- 3200
x"0e400",-- 3648
x"0b700",-- 2928
x"0eb00",-- 3760
x"0e400",-- 3648
x"0e200",-- 3616
x"11000",-- 4352
x"0fa00",-- 4000
x"0f800",-- 3968
x"0f400",-- 3904
x"0e900",-- 3728
x"0d800",-- 3456
x"0ce00",-- 3296
x"0b500",-- 2896
x"0a600",-- 2656
x"07b00",-- 1968
x"05c00",-- 1472
x"04400",-- 1088
x"01200",-- 288
x"ffd00",-- -48
x"fcc00",-- -832
x"fb200",-- -1248
x"f9500",-- -1712
x"f7c00",-- -2112
x"f6600",-- -2464
x"f3d00",-- -3120
x"f3000",-- -3328
x"f1c00",-- -3648
x"f1900",-- -3696
x"f0800",-- -3968
x"f0800",-- -3968
x"f0000",-- -4096
x"eff00",-- -4112
x"f0d00",-- -3888
x"f0d00",-- -3888
x"f1000",-- -3840
x"f2000",-- -3584
x"f3000",-- -3328
x"f3c00",-- -3136
x"f5600",-- -2720
x"f6500",-- -2480
x"f7400",-- -2240
x"f6800",-- -2432
x"f9200",-- -1760
x"f9100",-- -1776
x"fa300",-- -1488
x"fc600",-- -928
x"fbc00",-- -1088
x"fd500",-- -688
x"fd400",-- -704
x"ff400",-- -192
x"00300",-- 48
x"fe200",-- -480
x"01500",-- 336
x"03500",-- 848
x"ffb00",-- -80
x"04400",-- 1088
x"02c00",-- 704
x"03100",-- 784
x"05000",-- 1280
x"05100",-- 1296
x"06c00",-- 1728
x"06600",-- 1632
x"08d00",-- 2256
x"08400",-- 2112
x"0a100",-- 2576
x"0ac00",-- 2752
x"0bb00",-- 2992
x"0b600",-- 2912
x"0db00",-- 3504
x"0cb00",-- 3248
x"0ce00",-- 3296
x"0d000",-- 3328
x"0bf00",-- 3056
x"0f900",-- 3984
x"0c500",-- 3152
x"0dd00",-- 3536
x"0c700",-- 3184
x"0b800",-- 2944
x"0bd00",-- 3024
x"09200",-- 2336
x"09400",-- 2368
x"06b00",-- 1712
x"06000",-- 1536
x"03a00",-- 928
x"03700",-- 880
x"00800",-- 128
x"ff000",-- -256
x"fd200",-- -736
x"fb400",-- -1216
x"fa600",-- -1440
x"f8700",-- -1936
x"f8200",-- -2016
x"f5a00",-- -2656
x"f5800",-- -2688
x"f3e00",-- -3104
x"f4600",-- -2976
x"f3600",-- -3232
x"f2800",-- -3456
x"f3700",-- -3216
x"f2a00",-- -3424
x"f3c00",-- -3136
x"f2c00",-- -3392
x"f3c00",-- -3136
x"f3c00",-- -3136
x"f5500",-- -2736
x"f4d00",-- -2864
x"f7700",-- -2192
x"f5c00",-- -2624
x"f6d00",-- -2352
x"fa800",-- -1408
x"f5100",-- -2800
x"fb600",-- -1184
x"f9d00",-- -1584
x"fa300",-- -1488
x"fb300",-- -1232
x"fcb00",-- -848
x"fca00",-- -864
x"fcd00",-- -816
x"ff900",-- -112
x"fba00",-- -1120
x"02d00",-- 720
x"00000",-- 0
x"ffe00",-- -32
x"03500",-- 848
x"01200",-- 288
x"02f00",-- 752
x"05200",-- 1312
x"04a00",-- 1184
x"06700",-- 1648
x"05900",-- 1424
x"06400",-- 1600
x"07800",-- 1920
x"07200",-- 1824
x"0a800",-- 2688
x"08900",-- 2192
x"0a700",-- 2672
x"09600",-- 2400
x"0b600",-- 2912
x"0bb00",-- 2992
x"09700",-- 2416
x"0b700",-- 2928
x"0ac00",-- 2752
x"0b400",-- 2880
x"0a200",-- 2592
x"0c200",-- 3104
x"09500",-- 2384
x"0a300",-- 2608
x"0a100",-- 2576
x"07b00",-- 1968
x"08400",-- 2112
x"06600",-- 1632
x"06900",-- 1680
x"04f00",-- 1264
x"04f00",-- 1264
x"02300",-- 560
x"01100",-- 272
x"fe600",-- -416
x"fdc00",-- -576
x"fd500",-- -688
x"fc200",-- -992
x"fb700",-- -1168
x"f8e00",-- -1824
x"f8d00",-- -1840
x"f6600",-- -2464
x"f7b00",-- -2128
x"f5e00",-- -2592
x"f6900",-- -2416
x"f5800",-- -2688
x"f5d00",-- -2608
x"f5500",-- -2736
x"f4e00",-- -2848
x"f5c00",-- -2624
x"f3700",-- -3216
x"f6d00",-- -2352
x"f4a00",-- -2912
x"f8600",-- -1952
x"f4400",-- -3008
x"f8c00",-- -1856
x"f5d00",-- -2608
x"f7800",-- -2176
x"f9c00",-- -1600
x"f7000",-- -2304
x"fcb00",-- -848
x"f7500",-- -2224
x"fc900",-- -880
x"fa900",-- -1392
x"fd000",-- -768
x"fc700",-- -912
x"fde00",-- -544
x"fee00",-- -288
x"ff900",-- -112
x"00500",-- 80
x"01200",-- 288
x"00d00",-- 208
x"01a00",-- 416
x"03600",-- 864
x"01a00",-- 416
x"06100",-- 1552
x"03800",-- 896
x"04400",-- 1088
x"06e00",-- 1760
x"03c00",-- 960
x"06500",-- 1616
x"07500",-- 1872
x"05500",-- 1360
x"09300",-- 2352
x"07b00",-- 1968
x"07500",-- 1872
x"09f00",-- 2544
x"06a00",-- 1696
x"0b100",-- 2832
x"08900",-- 2192
x"09100",-- 2320
x"0a900",-- 2704
x"07700",-- 1904
x"0a900",-- 2704
x"09700",-- 2416
x"0a600",-- 2656
x"08200",-- 2080
x"09300",-- 2352
x"07200",-- 1824
x"07b00",-- 1968
x"06600",-- 1632
x"06400",-- 1600
x"05200",-- 1312
x"02800",-- 640
x"03a00",-- 928
x"00700",-- 112
x"00f00",-- 240
x"fe900",-- -368
x"fe500",-- -432
x"fc200",-- -992
x"fc300",-- -976
x"fb000",-- -1280
x"f9700",-- -1680
x"f9900",-- -1648
x"f7c00",-- -2112
x"f8400",-- -1984
x"f7100",-- -2288
x"f8200",-- -2016
x"f5900",-- -2672
x"f8000",-- -2048
x"f5a00",-- -2656
x"f6300",-- -2512
x"f6c00",-- -2368
x"f6600",-- -2464
x"f6400",-- -2496
x"f7500",-- -2224
x"f8900",-- -1904
x"f5e00",-- -2592
x"fb100",-- -1264
x"f5a00",-- -2656
x"fad00",-- -1328
x"f9a00",-- -1632
x"f7700",-- -2192
x"fdb00",-- -592
x"fa500",-- -1456
x"fb900",-- -1136
x"fb600",-- -1184
x"ffa00",-- -96
x"fb700",-- -1168
x"fe700",-- -400
x"00900",-- 144
x"fcd00",-- -816
x"02d00",-- 720
x"fdf00",-- -528
x"03200",-- 800
x"fed00",-- -304
x"03000",-- 768
x"01600",-- 352
x"01100",-- 272
x"06500",-- 1616
x"ffd00",-- -48
x"06b00",-- 1712
x"03300",-- 816
x"04000",-- 1024
x"07300",-- 1840
x"03f00",-- 1008
x"07200",-- 1824
x"06f00",-- 1776
x"06f00",-- 1776
x"08500",-- 2128
x"06c00",-- 1728
x"07400",-- 1856
x"09100",-- 2320
x"07500",-- 1872
x"09000",-- 2304
x"08600",-- 2144
x"08100",-- 2064
x"08f00",-- 2288
x"07e00",-- 2016
x"08d00",-- 2256
x"07900",-- 1936
x"08900",-- 2192
x"06500",-- 1616
x"07600",-- 1888
x"06b00",-- 1712
x"04900",-- 1168
x"04d00",-- 1232
x"03600",-- 864
x"03400",-- 832
x"01a00",-- 416
x"01300",-- 304
x"ff600",-- -160
x"ff700",-- -144
x"fd400",-- -704
x"fd500",-- -688
x"fc600",-- -928
x"f9a00",-- -1632
x"fbe00",-- -1056
x"f9300",-- -1744
x"f8700",-- -1936
x"f9c00",-- -1600
x"f8600",-- -1952
x"f7500",-- -2224
x"f8300",-- -2000
x"f7400",-- -2240
x"f7600",-- -2208
x"f8500",-- -1968
x"f6f00",-- -2320
x"f8e00",-- -1824
x"f6e00",-- -2336
x"f9800",-- -1664
x"f7800",-- -2176
x"f9000",-- -1792
x"fb200",-- -1248
x"f7300",-- -2256
x"fc200",-- -992
x"f9e00",-- -1568
x"f9d00",-- -1584
x"fcf00",-- -784
x"fa600",-- -1440
x"fc200",-- -992
x"fd200",-- -736
x"fbf00",-- -1040
x"ff300",-- -208
x"fc700",-- -912
x"fff00",-- -16
x"fdf00",-- -528
x"fe900",-- -368
x"03000",-- 768
x"fd800",-- -640
x"02200",-- 544
x"ffe00",-- -32
x"02d00",-- 720
x"00600",-- 96
x"02400",-- 576
x"03700",-- 880
x"02000",-- 512
x"04c00",-- 1216
x"01800",-- 384
x"08500",-- 2128
x"01500",-- 336
x"06900",-- 1680
x"06200",-- 1568
x"03e00",-- 992
x"08a00",-- 2208
x"04400",-- 1088
x"07d00",-- 2000
x"07100",-- 1808
x"07700",-- 1904
x"06500",-- 1616
x"09400",-- 2368
x"06100",-- 1552
x"07700",-- 1904
x"08c00",-- 2240
x"05700",-- 1392
x"08d00",-- 2256
x"07900",-- 1936
x"06b00",-- 1712
x"06e00",-- 1760
x"06400",-- 1600
x"05800",-- 1408
x"05400",-- 1344
x"03c00",-- 960
x"03700",-- 880
x"03300",-- 816
x"02900",-- 656
x"01a00",-- 416
x"fec00",-- -320
x"00b00",-- 176
x"fd100",-- -752
x"fe400",-- -448
x"fdd00",-- -560
x"fb400",-- -1216
x"fc300",-- -976
x"fb500",-- -1200
x"f9d00",-- -1584
x"fa200",-- -1504
x"fa800",-- -1408
x"f8800",-- -1920
x"fad00",-- -1328
x"f8200",-- -2016
x"f9f00",-- -1552
x"f9100",-- -1776
x"f9600",-- -1696
x"f8500",-- -1968
x"f9300",-- -1744
x"f9800",-- -1664
x"f9700",-- -1680
x"f9c00",-- -1600
x"f9800",-- -1664
x"fa800",-- -1408
x"f8a00",-- -1888
x"fb000",-- -1280
x"f9f00",-- -1552
x"fac00",-- -1344
x"fa900",-- -1392
x"fb200",-- -1248
x"fd300",-- -720
x"f9d00",-- -1584
x"fdf00",-- -528
x"fc900",-- -880
x"fcc00",-- -832
x"fea00",-- -352
x"fdb00",-- -592
x"ff800",-- -128
x"fd900",-- -624
x"01c00",-- 448
x"fda00",-- -608
x"01d00",-- 464
x"00500",-- 80
x"01b00",-- 432
x"00b00",-- 176
x"03c00",-- 960
x"03000",-- 768
x"02500",-- 592
x"03c00",-- 960
x"04600",-- 1120
x"04500",-- 1104
x"03c00",-- 960
x"06e00",-- 1760
x"04800",-- 1152
x"06500",-- 1616
x"04c00",-- 1216
x"06e00",-- 1760
x"04e00",-- 1248
x"05b00",-- 1456
x"08100",-- 2064
x"04800",-- 1152
x"07c00",-- 1984
x"06b00",-- 1712
x"06500",-- 1616
x"06900",-- 1680
x"06100",-- 1552
x"06000",-- 1536
x"04b00",-- 1200
x"07500",-- 1872
x"04d00",-- 1232
x"07b00",-- 1968
x"03200",-- 800
x"05400",-- 1344
x"03900",-- 912
x"04100",-- 1040
x"03900",-- 912
x"01f00",-- 496
x"02c00",-- 704
x"00400",-- 64
x"02700",-- 624
x"fed00",-- -304
x"ffb00",-- -80
x"fd300",-- -720
x"fe500",-- -432
x"fcd00",-- -816
x"fbe00",-- -1056
x"fe200",-- -480
x"fa100",-- -1520
x"fc000",-- -1024
x"fa900",-- -1392
x"f9e00",-- -1568
x"fae00",-- -1312
x"f9300",-- -1744
x"fa700",-- -1424
x"f9a00",-- -1632
x"fa500",-- -1456
x"f9c00",-- -1600
x"f9200",-- -1760
x"f9200",-- -1760
x"fa400",-- -1472
x"f9900",-- -1648
x"f8f00",-- -1808
x"fb600",-- -1184
x"fa500",-- -1456
x"f8400",-- -1984
x"fd600",-- -672
x"f8900",-- -1904
x"fb700",-- -1168
x"fb300",-- -1232
x"fa600",-- -1440
x"fd200",-- -736
x"fce00",-- -800
x"fd400",-- -704
x"fce00",-- -800
x"fe700",-- -400
x"fdf00",-- -528
x"fda00",-- -608
x"fed00",-- -304
x"01500",-- 336
x"ff400",-- -192
x"00600",-- 96
x"01e00",-- 480
x"ff700",-- -144
x"01700",-- 368
x"02500",-- 592
x"01e00",-- 480
x"01000",-- 256
x"05800",-- 1408
x"03f00",-- 1008
x"00900",-- 144
x"06000",-- 1536
x"01a00",-- 416
x"03b00",-- 944
x"05b00",-- 1456
x"02500",-- 592
x"05600",-- 1376
x"06100",-- 1552
x"03000",-- 768
x"06400",-- 1600
x"04500",-- 1104
x"03c00",-- 960
x"05900",-- 1424
x"05e00",-- 1504
x"05a00",-- 1440
x"07100",-- 1808
x"05100",-- 1296
x"04e00",-- 1248
x"05900",-- 1424
x"03100",-- 784
x"06e00",-- 1760
x"05200",-- 1312
x"05200",-- 1312
x"06b00",-- 1712
x"03200",-- 800
x"05700",-- 1392
x"03400",-- 832
x"02100",-- 528
x"03900",-- 912
x"01300",-- 304
x"02600",-- 608
x"01200",-- 288
x"00300",-- 48
x"ff500",-- -176
x"ff300",-- -208
x"fd100",-- -752
x"fe700",-- -400
x"fbb00",-- -1104
x"fd600",-- -672
x"fd500",-- -688
x"fa500",-- -1456
x"fd300",-- -720
x"fa300",-- -1488
x"fa000",-- -1536
x"fbc00",-- -1088
x"f9400",-- -1728
x"fae00",-- -1312
x"fba00",-- -1120
x"f9a00",-- -1632
x"f9f00",-- -1552
x"fac00",-- -1344
x"f8700",-- -1936
x"fae00",-- -1312
x"fbc00",-- -1088
x"f7500",-- -2224
x"fdb00",-- -592
x"fa300",-- -1488
x"fab00",-- -1360
x"faf00",-- -1296
x"fb500",-- -1200
x"faf00",-- -1296
x"fd300",-- -720
x"fc100",-- -1008
x"fbf00",-- -1040
x"fe500",-- -432
x"fa300",-- -1488
x"01200",-- 288
x"f9800",-- -1664
x"00500",-- 80
x"00000",-- 0
x"fd500",-- -688
x"00900",-- 144
x"fed00",-- -304
x"00d00",-- 208
x"00100",-- 16
x"01800",-- 384
x"ff600",-- -160
x"03700",-- 880
x"00400",-- 64
x"01300",-- 304
x"04b00",-- 1200
x"00000",-- 0
x"03a00",-- 928
x"02800",-- 640
x"03400",-- 832
x"03700",-- 880
x"02d00",-- 720
x"05b00",-- 1456
x"02f00",-- 752
x"03f00",-- 1008
x"04900",-- 1168
x"03600",-- 864
x"03800",-- 896
x"05600",-- 1376
x"03b00",-- 944
x"06b00",-- 1712
x"02500",-- 592
x"05900",-- 1424
x"04800",-- 1152
x"02b00",-- 688
x"07700",-- 1904
x"03700",-- 880
x"05300",-- 1328
x"04800",-- 1152
x"03800",-- 896
x"03900",-- 912
x"05b00",-- 1456
x"03800",-- 896
x"04100",-- 1040
x"03700",-- 880
x"03300",-- 816
x"03b00",-- 944
x"02500",-- 592
x"02700",-- 624
x"00800",-- 128
x"01c00",-- 448
x"fed00",-- -304
x"01400",-- 320
x"fe300",-- -464
x"fed00",-- -304
x"fec00",-- -320
x"fd100",-- -752
x"fde00",-- -544
x"fbd00",-- -1072
x"fcf00",-- -784
x"fb700",-- -1168
x"fc200",-- -992
x"fbb00",-- -1104
x"fc100",-- -1008
x"f9500",-- -1712
x"fb700",-- -1168
x"fab00",-- -1360
x"fbe00",-- -1056
x"f8f00",-- -1808
x"fd700",-- -656
x"f9d00",-- -1584
x"fa000",-- -1536
x"fd300",-- -720
x"f9500",-- -1712
x"fc500",-- -944
x"f9d00",-- -1584
x"fd100",-- -752
x"fa700",-- -1424
x"fcc00",-- -832
x"fb400",-- -1216
x"fbe00",-- -1056
x"fda00",-- -608
x"fa300",-- -1488
x"ffd00",-- -48
x"fb700",-- -1168
x"ffb00",-- -80
x"fbd00",-- -1072
x"fdb00",-- -592
x"ff500",-- -176
x"fd500",-- -688
x"00600",-- 96
x"fdc00",-- -576
x"01400",-- 320
x"fd200",-- -736
x"02400",-- 576
x"ff900",-- -112
x"00600",-- 96
x"01100",-- 272
x"01700",-- 368
x"01800",-- 384
x"00e00",-- 224
x"02100",-- 528
x"00e00",-- 224
x"03e00",-- 992
x"00d00",-- 208
x"04800",-- 1152
x"01f00",-- 496
x"03400",-- 832
x"03e00",-- 992
x"01600",-- 352
x"05f00",-- 1520
x"01700",-- 368
x"04700",-- 1136
x"03600",-- 864
x"04700",-- 1136
x"02800",-- 640
x"04200",-- 1056
x"06600",-- 1632
x"01900",-- 400
x"05f00",-- 1520
x"02a00",-- 672
x"06a00",-- 1696
x"02000",-- 512
x"05c00",-- 1472
x"03a00",-- 928
x"03900",-- 912
x"06400",-- 1600
x"01400",-- 320
x"06900",-- 1680
x"02300",-- 560
x"05200",-- 1312
x"02f00",-- 752
x"04500",-- 1104
x"03200",-- 800
x"00e00",-- 224
x"05300",-- 1328
x"fe000",-- -512
x"03f00",-- 1008
x"ff800",-- -128
x"ffa00",-- -96
x"01300",-- 304
x"fd900",-- -624
x"ff000",-- -256
x"fcd00",-- -816
x"fd800",-- -640
x"fc100",-- -1008
x"fef00",-- -272
x"fa600",-- -1440
x"fca00",-- -864
x"fcc00",-- -832
x"f8900",-- -1904
x"fc800",-- -896
x"fb500",-- -1200
x"faf00",-- -1296
x"fb500",-- -1200
x"fb500",-- -1200
x"f9300",-- -1744
x"fdb00",-- -592
x"f8c00",-- -1856
x"fc100",-- -1008
x"fcf00",-- -784
x"f9400",-- -1728
x"fe800",-- -384
x"f9100",-- -1776
x"fd600",-- -672
x"fb000",-- -1280
x"fb500",-- -1200
x"fe000",-- -512
x"fb500",-- -1200
x"fde00",-- -544
x"fe400",-- -448
x"fb100",-- -1264
x"fdd00",-- -560
x"ff300",-- -208
x"fb300",-- -1232
x"01100",-- 272
x"fe000",-- -512
x"fd900",-- -624
x"00800",-- 128
x"fdb00",-- -592
x"fff00",-- -16
x"00600",-- 96
x"fe400",-- -448
x"02f00",-- 752
x"00700",-- 112
x"fec00",-- -320
x"04e00",-- 1248
x"fe500",-- -432
x"01f00",-- 496
x"03000",-- 768
x"01000",-- 256
x"02200",-- 544
x"02f00",-- 752
x"02e00",-- 736
x"03300",-- 816
x"01a00",-- 416
x"03500",-- 848
x"04500",-- 1104
x"02c00",-- 704
x"04600",-- 1120
x"05b00",-- 1456
x"00f00",-- 240
x"05e00",-- 1504
x"03700",-- 880
x"02c00",-- 704
x"06800",-- 1664
x"03900",-- 912
x"05800",-- 1408
x"02800",-- 640
x"06a00",-- 1696
x"04800",-- 1152
x"04200",-- 1056
x"07000",-- 1792
x"02c00",-- 704
x"06100",-- 1552
x"05200",-- 1312
x"06200",-- 1568
x"04900",-- 1168
x"04600",-- 1120
x"06800",-- 1664
x"01c00",-- 448
x"04f00",-- 1264
x"03200",-- 800
x"04000",-- 1024
x"00d00",-- 208
x"01c00",-- 448
x"01c00",-- 448
x"fe200",-- -480
x"01300",-- 304
x"fc800",-- -896
x"ff500",-- -176
x"fc500",-- -944
x"fcd00",-- -816
x"fce00",-- -800
x"fb500",-- -1200
x"fc100",-- -1008
x"fad00",-- -1328
x"fc600",-- -928
x"f9d00",-- -1584
x"fbb00",-- -1104
x"fa500",-- -1456
x"fa800",-- -1408
x"f9900",-- -1648
x"fcb00",-- -848
x"f9600",-- -1696
x"fae00",-- -1312
x"fce00",-- -800
x"f9600",-- -1696
x"fc900",-- -880
x"faa00",-- -1376
x"fbf00",-- -1040
x"fac00",-- -1344
x"fc700",-- -912
x"fb600",-- -1184
x"fbf00",-- -1040
x"fdf00",-- -528
x"fab00",-- -1360
x"fd900",-- -624
x"fb300",-- -1232
x"fd700",-- -656
x"fe800",-- -384
x"fbf00",-- -1040
x"fc100",-- -1008
x"ffa00",-- -96
x"fca00",-- -864
x"ff500",-- -176
x"fdc00",-- -576
x"fd700",-- -656
x"01d00",-- 464
x"fcc00",-- -832
x"01c00",-- 448
x"fca00",-- -864
x"05500",-- 1360
x"fc800",-- -896
x"01600",-- 352
x"01c00",-- 448
x"fe600",-- -416
x"04300",-- 1072
x"00f00",-- 240
x"03a00",-- 928
x"ffd00",-- -48
x"05300",-- 1328
x"ff500",-- -176
x"03400",-- 832
x"04900",-- 1168
x"03600",-- 864
x"03100",-- 784
x"03d00",-- 976
x"05800",-- 1408
x"02100",-- 528
x"03500",-- 848
x"05c00",-- 1472
x"04d00",-- 1232
x"03f00",-- 1008
x"06f00",-- 1776
x"03a00",-- 928
x"05900",-- 1424
x"06100",-- 1552
x"04900",-- 1168
x"08600",-- 2144
x"03d00",-- 976
x"06f00",-- 1776
x"04c00",-- 1216
x"06800",-- 1664
x"08000",-- 2048
x"03a00",-- 928
x"07700",-- 1904
x"04600",-- 1120
x"05600",-- 1376
x"05600",-- 1376
x"05f00",-- 1520
x"01500",-- 336
x"03e00",-- 992
x"02200",-- 544
x"00a00",-- 160
x"02f00",-- 752
x"fea00",-- -352
x"00400",-- 64
x"fcf00",-- -784
x"fc500",-- -944
x"fcf00",-- -784
x"fc300",-- -976
x"fac00",-- -1344
x"fae00",-- -1312
x"fab00",-- -1360
x"faa00",-- -1376
x"f9100",-- -1776
x"f9b00",-- -1616
x"f9b00",-- -1616
x"f9800",-- -1664
x"fb300",-- -1232
x"f8e00",-- -1824
x"fac00",-- -1344
x"f9400",-- -1728
x"f9a00",-- -1632
x"fb100",-- -1264
x"fb800",-- -1152
x"fa300",-- -1488
x"fb100",-- -1264
x"fc100",-- -1008
x"fa700",-- -1424
x"fd000",-- -768
x"fae00",-- -1312
x"fac00",-- -1344
x"fda00",-- -608
x"fcb00",-- -848
x"f8e00",-- -1824
x"00d00",-- 208
x"fbb00",-- -1104
x"f8f00",-- -1808
x"fe900",-- -368
x"fd800",-- -640
x"fba00",-- -1120
x"fec00",-- -320
x"ffb00",-- -80
x"fc000",-- -1024
x"fdd00",-- -560
x"ff900",-- -112
x"fec00",-- -320
x"fe300",-- -464
x"01e00",-- 480
x"fe700",-- -400
x"03200",-- 800
x"fd100",-- -752
x"04200",-- 1056
x"00000",-- 0
x"ff100",-- -240
x"08400",-- 2112
x"fd000",-- -768
x"04900",-- 1168
x"02c00",-- 704
x"fe700",-- -400
x"05900",-- 1424
x"04100",-- 1040
x"ff300",-- -208
x"05f00",-- 1520
x"03700",-- 880
x"01600",-- 352
x"05a00",-- 1440
x"05100",-- 1296
x"03800",-- 896
x"05600",-- 1376
x"04000",-- 1024
x"07400",-- 1856
x"02500",-- 592
x"09300",-- 2352
x"06700",-- 1648
x"02b00",-- 688
x"0e200",-- 3616
x"02500",-- 592
x"07600",-- 1888
x"0ac00",-- 2752
x"05600",-- 1376
x"07d00",-- 2000
x"0b300",-- 2864
x"06900",-- 1680
x"07000",-- 1792
x"09100",-- 2320
x"04c00",-- 1216
x"08600",-- 2144
x"03f00",-- 1008
x"04900",-- 1168
x"03b00",-- 944
x"ffe00",-- -32
x"02c00",-- 704
x"feb00",-- -336
x"fed00",-- -304
x"fd300",-- -720
x"fa900",-- -1392
x"fb600",-- -1184
x"faf00",-- -1296
x"f8d00",-- -1840
x"f9000",-- -1792
x"f7e00",-- -2080
x"f7b00",-- -2128
x"f8100",-- -2032
x"f6800",-- -2432
x"f9e00",-- -1568
x"f6e00",-- -2336
x"f8700",-- -1936
x"f8800",-- -1920
x"f7f00",-- -2064
x"fa400",-- -1472
x"f8600",-- -1952
x"fb500",-- -1200
x"f9d00",-- -1584
x"faa00",-- -1376
x"fc100",-- -1008
x"fab00",-- -1360
x"fb700",-- -1168
x"fc000",-- -1024
x"fab00",-- -1360
x"fdf00",-- -528
x"fb300",-- -1232
x"fe200",-- -480
x"fc900",-- -880
x"f8600",-- -1952
x"ffd00",-- -48
x"fbb00",-- -1104
x"fbe00",-- -1056
x"fd700",-- -656
x"fd300",-- -720
x"fd500",-- -688
x"fbc00",-- -1088
x"fce00",-- -800
x"ffd00",-- -48
x"fab00",-- -1360
x"ff600",-- -160
x"00300",-- 48
x"fd900",-- -624
x"01e00",-- 480
x"fde00",-- -544
x"fe000",-- -512
x"03500",-- 848
x"fdd00",-- -560
x"00300",-- 48
x"03800",-- 896
x"01f00",-- 496
x"ff800",-- -128
x"05f00",-- 1520
x"fdf00",-- -528
x"03f00",-- 1008
x"05a00",-- 1440
x"fe800",-- -384
x"0b800",-- 2944
x"ffe00",-- -32
x"06000",-- 1536
x"04d00",-- 1232
x"01b00",-- 432
x"09200",-- 2336
x"03400",-- 832
x"08600",-- 2144
x"06c00",-- 1728
x"05600",-- 1376
x"0b900",-- 2960
x"04700",-- 1136
x"07d00",-- 2000
x"0ad00",-- 2768
x"0a900",-- 2704
x"08e00",-- 2272
x"08100",-- 2064
x"09b00",-- 2480
x"08c00",-- 2240
x"0a800",-- 2688
x"09200",-- 2336
x"0b400",-- 2880
x"0a200",-- 2592
x"04e00",-- 1248
x"0ab00",-- 2736
x"04f00",-- 1264
x"05800",-- 1408
x"05300",-- 1328
x"ffe00",-- -32
x"04300",-- 1072
x"fee00",-- -288
x"fdf00",-- -528
x"fc400",-- -960
x"f9f00",-- -1552
x"f9700",-- -1680
x"f8900",-- -1904
x"f8900",-- -1904
x"f7700",-- -2192
x"f5000",-- -2816
x"f5500",-- -2736
x"f5c00",-- -2624
x"f4c00",-- -2880
x"f6600",-- -2464
x"f6100",-- -2544
x"f6c00",-- -2368
x"f6700",-- -2448
x"f7500",-- -2224
x"f8200",-- -2016
x"f8400",-- -1984
x"f8a00",-- -1888
x"fa200",-- -1504
x"fb200",-- -1248
x"fac00",-- -1344
x"fbc00",-- -1088
x"fbb00",-- -1104
x"fb900",-- -1136
x"fd200",-- -736
x"fcd00",-- -816
x"fc700",-- -912
x"fdc00",-- -576
x"fc600",-- -928
x"fb600",-- -1184
x"feb00",-- -336
x"fda00",-- -608
x"fc700",-- -912
x"fd000",-- -768
x"fb500",-- -1200
x"fe600",-- -416
x"fbb00",-- -1104
x"fcf00",-- -784
x"fcd00",-- -816
x"fab00",-- -1360
x"fde00",-- -544
x"fcd00",-- -816
x"fe400",-- -448
x"fe400",-- -448
x"fdf00",-- -528
x"00200",-- 32
x"fd200",-- -736
x"00e00",-- 224
x"01600",-- 352
x"00500",-- 80
x"01400",-- 320
x"01a00",-- 416
x"02f00",-- 752
x"00700",-- 112
x"04e00",-- 1248
x"04b00",-- 1200
x"02000",-- 512
x"08300",-- 2096
x"06800",-- 1664
x"00a00",-- 160
x"09b00",-- 2480
x"05300",-- 1328
x"07300",-- 1840
x"0a500",-- 2640
x"05f00",-- 1520
x"0a700",-- 2672
x"06500",-- 1616
x"0ad00",-- 2768
x"0c000",-- 3072
x"0b100",-- 2832
x"0cd00",-- 3280
x"0c000",-- 3072
x"0a000",-- 2560
x"08c00",-- 2240
x"0ec00",-- 3776
x"0c800",-- 3200
x"0d100",-- 3344
x"0c700",-- 3184
x"09e00",-- 2528
x"0a200",-- 2592
x"08400",-- 2112
x"0a600",-- 2656
x"06d00",-- 1744
x"04d00",-- 1232
x"04200",-- 1056
x"fff00",-- -16
x"ff900",-- -112
x"fda00",-- -608
x"fa500",-- -1456
x"fa100",-- -1520
x"f8100",-- -2032
x"f5d00",-- -2608
x"f6600",-- -2464
x"f2e00",-- -3360
x"f3600",-- -3232
x"f2500",-- -3504
x"f2e00",-- -3360
x"f3c00",-- -3136
x"f3000",-- -3328
x"f2500",-- -3504
x"f3000",-- -3328
x"f3e00",-- -3104
x"f4700",-- -2960
x"f6600",-- -2464
x"f5f00",-- -2576
x"f7900",-- -2160
x"f7b00",-- -2128
x"f9a00",-- -1632
x"fa700",-- -1424
x"fad00",-- -1328
x"fb500",-- -1200
x"fbb00",-- -1104
x"fc500",-- -944
x"fd700",-- -656
x"fe700",-- -400
x"fde00",-- -544
x"fe100",-- -496
x"fe900",-- -368
x"fe700",-- -400
x"00500",-- 80
x"ff100",-- -240
x"ff200",-- -224
x"fdb00",-- -592
x"ff500",-- -176
x"fed00",-- -304
x"fd600",-- -672
x"ff900",-- -112
x"fdd00",-- -560
x"feb00",-- -336
x"ff000",-- -256
x"fd000",-- -768
x"fd900",-- -624
x"fef00",-- -272
x"fe900",-- -368
x"ff000",-- -256
x"ff900",-- -112
x"fd900",-- -624
x"ff100",-- -240
x"ffb00",-- -80
x"00800",-- 128
x"02400",-- 576
x"ffc00",-- -64
x"02600",-- 608
x"00d00",-- 208
x"03200",-- 800
x"04b00",-- 1200
x"04d00",-- 1232
x"05400",-- 1344
x"05c00",-- 1472
x"07600",-- 1888
x"06f00",-- 1776
x"08500",-- 2128
x"08700",-- 2160
x"09c00",-- 2496
x"0a200",-- 2592
x"0a800",-- 2688
x"0cf00",-- 3312
x"0c300",-- 3120
x"0cb00",-- 3248
x"10400",-- 4160
x"0e800",-- 3712
x"09600",-- 2400
x"0c500",-- 3152
x"0ec00",-- 3776
x"0ed00",-- 3792
x"0f400",-- 3904
x"0d900",-- 3472
x"0ad00",-- 2768
x"08600",-- 2144
x"09300",-- 2352
x"0a300",-- 2608
x"09a00",-- 2464
x"04f00",-- 1264
x"01b00",-- 432
x"ff900",-- -112
x"fd700",-- -656
x"fc700",-- -912
x"fae00",-- -1312
x"f8300",-- -2000
x"f6200",-- -2528
x"f3c00",-- -3136
x"f2a00",-- -3424
x"f1f00",-- -3600
x"efc00",-- -4160
x"f0200",-- -4064
x"f1f00",-- -3600
x"f1b00",-- -3664
x"f1600",-- -3744
x"f0000",-- -4096
x"f0b00",-- -3920
x"f2000",-- -3584
x"f4000",-- -3072
x"f6100",-- -2544
x"f6500",-- -2480
x"f5a00",-- -2656
x"f5900",-- -2672
x"f8700",-- -1936
x"fa400",-- -1472
x"fb000",-- -1280
x"fbe00",-- -1056
x"fc500",-- -944
x"fc600",-- -928
x"fce00",-- -800
x"fde00",-- -544
x"fe500",-- -432
x"ff200",-- -224
x"00000",-- 0
x"00900",-- 144
x"ff400",-- -192
x"fd700",-- -656
x"fe300",-- -464
x"fff00",-- -16
x"01200",-- 288
x"01100",-- 272
x"ff400",-- -192
x"fca00",-- -864
x"fdd00",-- -560
x"ff000",-- -256
x"00800",-- 128
x"00000",-- 0
x"fe200",-- -480
x"fe900",-- -368
x"fe900",-- -368
x"fe300",-- -464
x"ffc00",-- -64
x"ffe00",-- -32
x"ff300",-- -208
x"01100",-- 272
x"01200",-- 288
x"00100",-- 16
x"00a00",-- 160
x"02000",-- 512
x"03000",-- 768
x"04600",-- 1120
x"05b00",-- 1456
x"04000",-- 1024
x"05500",-- 1360
x"06500",-- 1616
x"06e00",-- 1760
x"09900",-- 2448
x"0a500",-- 2640
x"09600",-- 2400
x"09d00",-- 2512
x"0c400",-- 3136
x"0dd00",-- 3536
x"0ff00",-- 4080
x"10400",-- 4160
x"0f700",-- 3952
x"0cb00",-- 3248
x"0c000",-- 3072
x"0e800",-- 3712
x"11a00",-- 4512
x"12f00",-- 4848
x"0f200",-- 3872
x"0d600",-- 3424
x"0ae00",-- 2784
x"09b00",-- 2480
x"0d000",-- 3328
x"0b100",-- 2832
x"07700",-- 1904
x"03900",-- 912
x"ff400",-- -192
x"fe900",-- -368
x"fc700",-- -912
x"fac00",-- -1344
x"f8c00",-- -1856
x"f6100",-- -2544
x"f3500",-- -3248
x"f1000",-- -3840
x"f0600",-- -4000
x"ef100",-- -4336
x"eec00",-- -4416
x"f0500",-- -4016
x"f0b00",-- -3920
x"ef100",-- -4336
x"edd00",-- -4656
x"ee500",-- -4528
x"f0500",-- -4016
x"f2800",-- -3456
x"f4400",-- -3008
x"f4600",-- -2976
x"f3600",-- -3232
x"f3c00",-- -3136
x"f6c00",-- -2368
x"f9c00",-- -1600
x"fa800",-- -1408
x"fab00",-- -1360
x"fb300",-- -1232
x"fb200",-- -1248
x"fb700",-- -1168
x"fdd00",-- -560
x"ff200",-- -224
x"00100",-- 16
x"fff00",-- -16
x"ff800",-- -128
x"ffc00",-- -64
x"ff700",-- -144
x"00f00",-- 240
x"02400",-- 576
x"02400",-- 576
x"01200",-- 288
x"00900",-- 144
x"fed00",-- -304
x"ff000",-- -256
x"01c00",-- 448
x"01c00",-- 448
x"02500",-- 592
x"ff500",-- -176
x"fd300",-- -720
x"ff600",-- -160
x"00a00",-- 160
x"00b00",-- 176
x"01400",-- 320
x"fef00",-- -272
x"fd500",-- -688
x"ff000",-- -256
x"00100",-- 16
x"01400",-- 320
x"01600",-- 352
x"00f00",-- 240
x"00800",-- 128
x"02100",-- 528
x"02900",-- 656
x"03a00",-- 928
x"06200",-- 1568
x"05400",-- 1344
x"07200",-- 1824
x"07200",-- 1824
x"07a00",-- 1952
x"0a400",-- 2624
x"0ac00",-- 2752
x"0d300",-- 3376
x"0e700",-- 3696
x"0d600",-- 3424
x"0fc00",-- 4032
x"10300",-- 4144
x"0cd00",-- 3280
x"0dd00",-- 3536
x"10500",-- 4176
x"11c00",-- 4544
x"12600",-- 4704
x"10300",-- 4144
x"0cf00",-- 3312
x"0bd00",-- 3024
x"0b800",-- 2944
x"0ce00",-- 3296
x"0c000",-- 3072
x"07700",-- 1904
x"01500",-- 336
x"fec00",-- -320
x"fef00",-- -272
x"fdb00",-- -592
x"fc300",-- -976
x"f8900",-- -1904
x"f4900",-- -2928
x"f1800",-- -3712
x"f1300",-- -3792
x"f1b00",-- -3664
x"f0a00",-- -3936
x"ef200",-- -4320
x"ef500",-- -4272
x"ef000",-- -4352
x"ee000",-- -4608
x"ee700",-- -4496
x"ef600",-- -4256
x"f1300",-- -3792
x"f2a00",-- -3424
x"f3900",-- -3184
x"f3000",-- -3328
x"f3100",-- -3312
x"f4300",-- -3024
x"f7300",-- -2256
x"fa800",-- -1408
x"fa700",-- -1424
x"f9600",-- -1696
x"f9400",-- -1728
x"fa700",-- -1424
x"fcb00",-- -848
x"fe600",-- -416
x"fea00",-- -352
x"fe600",-- -416
x"fe200",-- -480
x"00100",-- 16
x"00c00",-- 192
x"00800",-- 128
x"01200",-- 288
x"01400",-- 320
x"01f00",-- 496
x"02500",-- 592
x"01800",-- 384
x"00e00",-- 224
x"00800",-- 128
x"01300",-- 304
x"02d00",-- 720
x"02000",-- 512
x"fff00",-- -16
x"fee00",-- -288
x"ff300",-- -208
x"00600",-- 96
x"01600",-- 352
x"00e00",-- 224
x"ff100",-- -240
x"fe600",-- -416
x"ff100",-- -240
x"00100",-- 16
x"01300",-- 304
x"00800",-- 128
x"ffe00",-- -32
x"00f00",-- 240
x"01000",-- 256
x"02200",-- 544
x"03100",-- 784
x"03800",-- 896
x"05700",-- 1392
x"05c00",-- 1472
x"05f00",-- 1520
x"06900",-- 1680
x"07e00",-- 2016
x"09300",-- 2352
x"0c000",-- 3072
x"0d400",-- 3392
x"0c700",-- 3184
x"0e200",-- 3616
x"0fa00",-- 4000
x"0d800",-- 3456
x"0d900",-- 3472
x"0e900",-- 3728
x"0ee00",-- 3808
x"13400",-- 4928
x"12400",-- 4672
x"0e600",-- 3680
x"0c300",-- 3120
x"0a500",-- 2640
x"0c200",-- 3104
x"0dc00",-- 3520
x"0b600",-- 2912
x"05800",-- 1408
x"ff600",-- -160
x"fe300",-- -464
x"ffa00",-- -96
x"ff400",-- -192
x"fbd00",-- -1072
x"f6900",-- -2416
x"f2800",-- -3456
x"f0600",-- -4000
x"f1d00",-- -3632
x"f3500",-- -3248
x"f1700",-- -3728
x"ef700",-- -4240
x"ee300",-- -4560
x"ee200",-- -4576
x"eee00",-- -4384
x"ef700",-- -4240
x"f1300",-- -3792
x"f2900",-- -3440
x"f2600",-- -3488
x"f2500",-- -3504
x"f2600",-- -3488
x"f3300",-- -3280
x"f5c00",-- -2624
x"f8e00",-- -1824
x"fa900",-- -1392
x"f8b00",-- -1872
x"f7800",-- -2176
x"f9100",-- -1776
x"fba00",-- -1120
x"fe200",-- -480
x"ff500",-- -176
x"fdf00",-- -528
x"fba00",-- -1120
x"fd200",-- -736
x"00100",-- 16
x"02a00",-- 672
x"02c00",-- 704
x"00a00",-- 160
x"00500",-- 80
x"01000",-- 256
x"02800",-- 640
x"03b00",-- 944
x"03e00",-- 992
x"01400",-- 320
x"00900",-- 144
x"02800",-- 640
x"02300",-- 560
x"02c00",-- 704
x"01a00",-- 416
x"00500",-- 80
x"00e00",-- 224
x"00900",-- 144
x"00700",-- 112
x"00300",-- 48
x"fe900",-- -368
x"fec00",-- -320
x"fff00",-- -16
x"ffa00",-- -96
x"fe600",-- -416
x"fe600",-- -416
x"fea00",-- -352
x"ff400",-- -192
x"01000",-- 256
x"01000",-- 256
x"01100",-- 272
x"01500",-- 336
x"02500",-- 592
x"04f00",-- 1264
x"05a00",-- 1440
x"05a00",-- 1440
x"07500",-- 1872
x"08300",-- 2096
x"0a200",-- 2592
x"0b600",-- 2912
x"0be00",-- 3040
x"0e100",-- 3600
x"0f700",-- 3952
x"0f900",-- 3984
x"0f300",-- 3888
x"0d500",-- 3408
x"0ca00",-- 3232
x"10600",-- 4192
x"13600",-- 4960
x"12a00",-- 4768
x"0e300",-- 3632
x"09d00",-- 2512
x"0a800",-- 2688
x"0bf00",-- 3056
x"0cb00",-- 3248
x"0aa00",-- 2720
x"03900",-- 912
x"fe200",-- -480
x"fe200",-- -480
x"ff400",-- -192
x"fdf00",-- -528
x"fad00",-- -1328
x"f5c00",-- -2624
x"f1d00",-- -3632
x"f1b00",-- -3664
x"f2b00",-- -3408
x"f2d00",-- -3376
x"f1b00",-- -3664
x"eff00",-- -4112
x"eef00",-- -4368
x"efa00",-- -4192
x"efc00",-- -4160
x"f0500",-- -4016
x"f2200",-- -3552
x"f3200",-- -3296
x"f3700",-- -3216
x"f2f00",-- -3344
x"f2e00",-- -3360
x"f4300",-- -3024
x"f6e00",-- -2336
x"f9700",-- -1680
x"fa000",-- -1536
x"f8500",-- -1968
x"f7800",-- -2176
x"f9600",-- -1696
x"fce00",-- -800
x"fe400",-- -448
x"fe600",-- -416
x"fd800",-- -640
x"fc800",-- -896
x"fd900",-- -624
x"fff00",-- -16
x"02800",-- 640
x"02d00",-- 720
x"01b00",-- 432
x"00900",-- 144
x"00900",-- 144
x"01e00",-- 480
x"03400",-- 832
x"03b00",-- 944
x"03a00",-- 928
x"01a00",-- 416
x"00600",-- 96
x"00800",-- 128
x"01800",-- 384
x"03200",-- 800
x"02600",-- 608
x"00200",-- 32
x"fe200",-- -480
x"fd800",-- -640
x"ff900",-- -112
x"01100",-- 272
x"00f00",-- 240
x"fee00",-- -288
x"fd000",-- -768
x"fd400",-- -704
x"fea00",-- -352
x"00c00",-- 192
x"00f00",-- 240
x"ffc00",-- -64
x"ff300",-- -208
x"ff800",-- -128
x"01100",-- 272
x"03700",-- 880
x"05000",-- 1280
x"04e00",-- 1248
x"04a00",-- 1184
x"05a00",-- 1440
x"06f00",-- 1776
x"09500",-- 2384
x"0a600",-- 2656
x"0bd00",-- 3024
x"0d900",-- 3472
x"0cd00",-- 3280
x"0e400",-- 3648
x"10100",-- 4112
x"0e500",-- 3664
x"0dc00",-- 3520
x"0eb00",-- 3760
x"10a00",-- 4256
x"12500",-- 4688
x"10500",-- 4176
x"0ca00",-- 3232
x"0a300",-- 2608
x"0b500",-- 2896
x"0d800",-- 3456
x"0b600",-- 2912
x"06c00",-- 1728
x"01a00",-- 416
x"fed00",-- -304
x"ff200",-- -224
x"00000",-- 0
x"fdb00",-- -592
x"f7f00",-- -2064
x"f3f00",-- -3088
x"f2b00",-- -3408
x"f3600",-- -3232
x"f4300",-- -3024
x"f3000",-- -3328
x"f0e00",-- -3872
x"ef600",-- -4256
x"ef100",-- -4336
x"f0a00",-- -3936
x"f1600",-- -3744
x"f1600",-- -3744
x"f2200",-- -3552
x"f3200",-- -3296
x"f3300",-- -3280
x"f2800",-- -3456
x"f3500",-- -3248
x"f6000",-- -2560
x"f8000",-- -2048
x"f8f00",-- -1808
x"f8200",-- -2016
x"f7700",-- -2192
x"f8400",-- -1984
x"fb000",-- -1280
x"fe600",-- -416
x"fe700",-- -400
x"fc300",-- -976
x"fb800",-- -1152
x"fdb00",-- -592
x"00900",-- 144
x"02000",-- 512
x"00b00",-- 176
x"ffe00",-- -32
x"00d00",-- 208
x"02b00",-- 688
x"03b00",-- 944
x"02d00",-- 720
x"01d00",-- 464
x"02500",-- 592
x"03900",-- 912
x"03600",-- 864
x"02200",-- 544
x"00400",-- 64
x"ff900",-- -112
x"02a00",-- 672
x"03500",-- 848
x"00800",-- 128
x"fe100",-- -496
x"fcb00",-- -848
x"fee00",-- -288
x"01900",-- 400
x"00400",-- 64
x"fdd00",-- -560
x"fbb00",-- -1104
x"fc200",-- -992
x"ff400",-- -192
x"01300",-- 304
x"ffa00",-- -96
x"fd400",-- -704
x"fdb00",-- -592
x"ffa00",-- -96
x"01e00",-- 480
x"02f00",-- 752
x"02800",-- 640
x"02700",-- 624
x"03d00",-- 976
x"06500",-- 1616
x"08100",-- 2064
x"08200",-- 2080
x"08c00",-- 2240
x"0a000",-- 2560
x"0c600",-- 3168
x"0da00",-- 3488
x"0e500",-- 3664
x"0f200",-- 3872
x"0f300",-- 3888
x"10200",-- 4128
x"0e900",-- 3728
x"0e400",-- 3648
x"12500",-- 4688
x"13200",-- 4896
x"10f00",-- 4336
x"0cd00",-- 3280
x"0a600",-- 2656
x"0d100",-- 3344
x"0d300",-- 3376
x"0a300",-- 2608
x"07400",-- 1856
x"02400",-- 576
x"fe000",-- -512
x"fe500",-- -432
x"00d00",-- 208
x"fd400",-- -704
x"f6500",-- -2480
x"f4000",-- -3072
x"f2f00",-- -3344
x"f2f00",-- -3344
x"f3700",-- -3216
x"f3000",-- -3328
x"f1400",-- -3776
x"ee500",-- -4528
x"ee400",-- -4544
x"f1100",-- -3824
x"f1e00",-- -3616
x"f1500",-- -3760
x"f1f00",-- -3600
x"f3300",-- -3280
x"f2000",-- -3584
x"f1400",-- -3776
x"f4c00",-- -2880
x"f7500",-- -2224
x"f7a00",-- -2144
x"f7500",-- -2224
x"f7700",-- -2192
x"f7c00",-- -2112
x"f8700",-- -1936
x"fc500",-- -944
x"ff000",-- -256
x"fcc00",-- -832
x"fb500",-- -1200
x"fcd00",-- -816
x"fea00",-- -352
x"00b00",-- 176
x"02800",-- 640
x"02a00",-- 672
x"00300",-- 48
x"fe500",-- -432
x"01e00",-- 480
x"06400",-- 1600
x"06500",-- 1616
x"03400",-- 832
x"01200",-- 288
x"00a00",-- 160
x"01300",-- 304
x"05800",-- 1408
x"06400",-- 1600
x"01e00",-- 480
x"fd900",-- -624
x"fcc00",-- -832
x"00b00",-- 176
x"02800",-- 640
x"01400",-- 320
x"fec00",-- -320
x"fb500",-- -1200
x"fb000",-- -1280
x"fd800",-- -640
x"00800",-- 128
x"00500",-- 80
x"fcf00",-- -784
x"fc300",-- -976
x"fc900",-- -880
x"fe100",-- -496
x"00300",-- 48
x"01900",-- 400
x"01a00",-- 416
x"ff700",-- -144
x"ff900",-- -112
x"02400",-- 576
x"04d00",-- 1232
x"06f00",-- 1776
x"07400",-- 1856
x"06a00",-- 1696
x"06c00",-- 1728
x"08500",-- 2128
x"0c000",-- 3072
x"0e500",-- 3664
x"0e900",-- 3728
x"0ec00",-- 3776
x"0e000",-- 3584
x"0eb00",-- 3760
x"10700",-- 4208
x"0f600",-- 3936
x"0f000",-- 3840
x"12100",-- 4624
x"13300",-- 4912
x"10100",-- 4112
x"0ab00",-- 2736
x"0a400",-- 2624
x"0e400",-- 3648
x"0e300",-- 3632
x"09f00",-- 2544
x"05500",-- 1360
x"00400",-- 64
x"fdd00",-- -560
x"00000",-- 0
x"02000",-- 512
x"fcc00",-- -832
x"f4600",-- -2976
x"f1c00",-- -3648
x"f3b00",-- -3152
x"f5000",-- -2816
x"f3c00",-- -3136
x"f2900",-- -3440
x"f0600",-- -4000
x"ece00",-- -4896
x"ee300",-- -4560
x"f2900",-- -3440
x"f2d00",-- -3376
x"f0b00",-- -3920
x"f1500",-- -3760
x"f2d00",-- -3376
x"f1800",-- -3712
x"f1a00",-- -3680
x"f5a00",-- -2656
x"f8600",-- -1952
x"f7700",-- -2192
x"f6200",-- -2528
x"f6e00",-- -2336
x"f8400",-- -1984
x"f9b00",-- -1616
x"fda00",-- -608
x"ff400",-- -192
x"fbb00",-- -1104
x"fa000",-- -1536
x"fdc00",-- -576
x"01400",-- 320
x"01f00",-- 496
x"02100",-- 528
x"01800",-- 384
x"00000",-- 0
x"ff700",-- -144
x"03700",-- 880
x"07600",-- 1888
x"05500",-- 1360
x"02500",-- 592
x"01500",-- 336
x"02200",-- 544
x"03b00",-- 944
x"04f00",-- 1264
x"05000",-- 1280
x"01a00",-- 416
x"fd500",-- -688
x"fca00",-- -864
x"01c00",-- 448
x"03600",-- 864
x"00000",-- 0
x"fd100",-- -752
x"fa100",-- -1520
x"fab00",-- -1360
x"feb00",-- -336
x"00700",-- 112
x"fe700",-- -400
x"fa600",-- -1440
x"f9300",-- -1744
x"fc100",-- -1008
x"ff600",-- -160
x"ffc00",-- -64
x"fe200",-- -480
x"fdc00",-- -576
x"fd300",-- -720
x"fec00",-- -320
x"02b00",-- 688
x"04700",-- 1136
x"04200",-- 1056
x"03e00",-- 992
x"04800",-- 1152
x"06900",-- 1680
x"08f00",-- 2288
x"0b900",-- 2960
x"0c100",-- 3088
x"0bb00",-- 2992
x"0c400",-- 3136
x"0e500",-- 3664
x"10c00",-- 4288
x"11700",-- 4464
x"12200",-- 4640
x"10d00",-- 4304
x"0bd00",-- 3024
x"0e300",-- 3632
x"15700",-- 5488
x"15500",-- 5456
x"0fe00",-- 4064
x"08700",-- 2160
x"09500",-- 2384
x"0d800",-- 3456
x"0bf00",-- 3056
x"09c00",-- 2496
x"05200",-- 1312
x"fdd00",-- -560
x"faf00",-- -1296
x"fea00",-- -352
x"00a00",-- 160
x"f9900",-- -1648
x"f3600",-- -3232
x"f2e00",-- -3360
x"f1c00",-- -3648
x"f1200",-- -3808
x"f1b00",-- -3664
x"f3100",-- -3312
x"f0600",-- -4000
x"ebe00",-- -5152
x"ede00",-- -4640
x"f0c00",-- -3904
x"f0200",-- -4064
x"f1300",-- -3792
x"f3c00",-- -3136
x"f2b00",-- -3408
x"eef00",-- -4368
x"f1000",-- -3840
x"f7400",-- -2240
x"f9000",-- -1792
x"f7a00",-- -2144
x"f7000",-- -2304
x"f7600",-- -2208
x"f7800",-- -2176
x"fac00",-- -1344
x"00600",-- 96
x"ff800",-- -128
x"fb500",-- -1200
x"fbe00",-- -1056
x"ff900",-- -112
x"01b00",-- 432
x"02600",-- 608
x"03700",-- 880
x"02c00",-- 704
x"00e00",-- 224
x"02100",-- 528
x"05000",-- 1280
x"04500",-- 1104
x"03700",-- 880
x"05400",-- 1344
x"05400",-- 1344
x"02a00",-- 672
x"00300",-- 48
x"02200",-- 544
x"03c00",-- 960
x"02600",-- 608
x"00b00",-- 176
x"fe900",-- -368
x"fd400",-- -704
x"fbb00",-- -1104
x"fe800",-- -384
x"00f00",-- 240
x"fc100",-- -1008
x"f9500",-- -1712
x"fa300",-- -1488
x"fb000",-- -1280
x"fca00",-- -864
x"fd500",-- -688
x"fd200",-- -736
x"fb200",-- -1248
x"fa800",-- -1408
x"fd600",-- -672
x"ffb00",-- -80
x"00700",-- 112
x"ff900",-- -112
x"00800",-- 128
x"02200",-- 544
x"02700",-- 624
x"04d00",-- 1232
x"07800",-- 1920
x"07c00",-- 1984
x"07b00",-- 1968
x"09000",-- 2304
x"0bb00",-- 2992
x"0c300",-- 3120
x"0cf00",-- 3312
x"0f400",-- 3904
x"10500",-- 4176
x"10900",-- 4240
x"10c00",-- 4288
x"11a00",-- 4512
x"12600",-- 4704
x"0e800",-- 3712
x"0d100",-- 3344
x"13e00",-- 5088
x"15400",-- 5440
x"10000",-- 4096
x"08f00",-- 2288
x"08b00",-- 2224
x"0d300",-- 3376
x"0c100",-- 3088
x"09900",-- 2448
x"04e00",-- 1248
x"fd500",-- -688
x"fa800",-- -1408
x"fdd00",-- -560
x"00a00",-- 160
x"fa900",-- -1392
x"f1800",-- -3712
x"f0500",-- -4016
x"f1b00",-- -3664
x"f1900",-- -3696
x"f0e00",-- -3872
x"f1400",-- -3776
x"eef00",-- -4368
x"ea300",-- -5584
x"ecc00",-- -4928
x"f1800",-- -3712
x"f0300",-- -4048
x"eef00",-- -4368
x"f1800",-- -3712
x"f2d00",-- -3376
x"f0400",-- -4032
x"f0e00",-- -3872
x"f6700",-- -2448
x"f8b00",-- -1872
x"f7b00",-- -2128
x"f7900",-- -2160
x"f8d00",-- -1840
x"f9300",-- -1744
x"faf00",-- -1296
x"00100",-- 16
x"01600",-- 352
x"fd400",-- -704
x"fc900",-- -880
x"00900",-- 144
x"03d00",-- 976
x"03800",-- 896
x"03400",-- 832
x"04800",-- 1152
x"01a00",-- 416
x"01b00",-- 432
x"06000",-- 1536
x"06e00",-- 1760
x"05200",-- 1312
x"03100",-- 784
x"03200",-- 800
x"03c00",-- 960
x"02600",-- 608
x"02900",-- 656
x"03200",-- 800
x"01b00",-- 432
x"fe200",-- -480
x"fc300",-- -976
x"ff200",-- -224
x"fe100",-- -496
x"fdf00",-- -528
x"fe000",-- -512
x"f9700",-- -1680
x"f8b00",-- -1872
x"fa600",-- -1440
x"fd500",-- -688
x"fd900",-- -624
x"fa400",-- -1472
x"f9100",-- -1776
x"f9d00",-- -1584
x"fc600",-- -928
x"fea00",-- -352
x"ff000",-- -256
x"fe900",-- -368
x"fcd00",-- -816
x"fe800",-- -384
x"02800",-- 640
x"04d00",-- 1232
x"05400",-- 1344
x"05100",-- 1296
x"06500",-- 1616
x"07000",-- 1792
x"09100",-- 2320
x"0ca00",-- 3232
x"0d600",-- 3424
x"0ca00",-- 3232
x"0d100",-- 3344
x"0e500",-- 3664
x"10400",-- 4160
x"12600",-- 4704
x"12800",-- 4736
x"12f00",-- 4848
x"11d00",-- 4560
x"10300",-- 4144
x"0d100",-- 3344
x"0eb00",-- 3760
x"15c00",-- 5568
x"13c00",-- 5056
x"0dc00",-- 3520
x"06e00",-- 1760
x"06200",-- 1568
x"0bd00",-- 3024
x"0b700",-- 2928
x"07e00",-- 2016
x"01900",-- 400
x"f9400",-- -1728
x"f7900",-- -2160
x"fbc00",-- -1088
x"fee00",-- -288
x"f8200",-- -2016
x"eed00",-- -4400
x"edd00",-- -4656
x"ede00",-- -4640
x"eee00",-- -4384
x"f1000",-- -3840
x"f0a00",-- -3936
x"ec600",-- -5024
x"e8c00",-- -5952
x"ec200",-- -5088
x"f0000",-- -4096
x"f0100",-- -4080
x"f0c00",-- -3904
x"f2600",-- -3488
x"f2900",-- -3440
x"f0c00",-- -3904
x"f2300",-- -3536
x"f8400",-- -1984
x"faf00",-- -1296
x"fa500",-- -1456
x"fa600",-- -1440
x"fa700",-- -1424
x"fa500",-- -1456
x"fd800",-- -640
x"03c00",-- 960
x"04400",-- 1088
x"ffd00",-- -48
x"ff100",-- -240
x"01700",-- 368
x"04000",-- 1024
x"06700",-- 1648
x"07100",-- 1808
x"05800",-- 1408
x"02500",-- 592
x"02500",-- 592
x"04000",-- 1024
x"06100",-- 1552
x"07b00",-- 1968
x"04500",-- 1104
x"02a00",-- 672
x"fff00",-- -16
x"fdf00",-- -528
x"02c00",-- 704
x"04500",-- 1104
x"00400",-- 64
x"fae00",-- -1312
x"f8e00",-- -1824
x"fa600",-- -1440
x"fd100",-- -752
x"ff100",-- -240
x"fb700",-- -1168
x"f7200",-- -2272
x"f6600",-- -2464
x"f8200",-- -2016
x"fc700",-- -912
x"fd000",-- -768
x"fa600",-- -1440
x"f9500",-- -1712
x"f9b00",-- -1616
x"fc500",-- -944
x"fec00",-- -320
x"00900",-- 144
x"00c00",-- 192
x"ffc00",-- -64
x"01300",-- 304
x"03500",-- 848
x"05900",-- 1424
x"07e00",-- 2016
x"09600",-- 2400
x"09e00",-- 2528
x"09200",-- 2336
x"0aa00",-- 2720
x"0d400",-- 3392
x"0eb00",-- 3760
x"10b00",-- 4272
x"0f600",-- 3936
x"0ef00",-- 3824
x"11100",-- 4368
x"11e00",-- 4576
x"13700",-- 4976
x"14600",-- 5216
x"12800",-- 4736
x"10f00",-- 4336
x"0d400",-- 3392
x"0be00",-- 3040
x"12b00",-- 4784
x"13e00",-- 5088
x"0fb00",-- 4016
x"07700",-- 1904
x"03600",-- 864
x"07a00",-- 1952
x"08400",-- 2112
x"07300",-- 1840
x"02f00",-- 752
x"f9900",-- -1648
x"f4600",-- -2976
x"f6000",-- -2560
x"fa700",-- -1424
x"f8800",-- -1920
x"f0500",-- -4016
x"ec300",-- -5072
x"ea800",-- -5504
x"eaf00",-- -5392
x"ed700",-- -4752
x"ef800",-- -4224
x"ee000",-- -4608
x"e9300",-- -5840
x"e9d00",-- -5680
x"edc00",-- -4672
x"ef400",-- -4288
x"f0700",-- -3984
x"f3700",-- -3216
x"f4f00",-- -2832
x"f2f00",-- -3344
x"f2800",-- -3456
x"f7200",-- -2272
x"fb400",-- -1216
x"fd100",-- -752
x"fe600",-- -416
x"fe500",-- -432
x"fc600",-- -928
x"fcf00",-- -784
x"02e00",-- 736
x"07000",-- 1792
x"05900",-- 1424
x"02f00",-- 752
x"02200",-- 544
x"02600",-- 608
x"04d00",-- 1232
x"08000",-- 2048
x"08f00",-- 2288
x"05200",-- 1312
x"00900",-- 144
x"01f00",-- 496
x"05500",-- 1360
x"05f00",-- 1520
x"04600",-- 1120
x"01f00",-- 496
x"ff400",-- -192
x"fd200",-- -736
x"ff100",-- -240
x"00900",-- 144
x"fdb00",-- -592
x"fbf00",-- -1040
x"f9a00",-- -1632
x"fa800",-- -1408
x"fa400",-- -1472
x"f8500",-- -1968
x"fb600",-- -1184
x"f9d00",-- -1584
x"f8c00",-- -1856
x"f9700",-- -1680
x"f8c00",-- -1856
x"f9f00",-- -1552
x"fad00",-- -1328
x"fd400",-- -704
x"fe300",-- -464
x"fc800",-- -896
x"fca00",-- -864
x"feb00",-- -336
x"02600",-- 608
x"03f00",-- 1008
x"03e00",-- 992
x"04b00",-- 1200
x"04900",-- 1168
x"06c00",-- 1728
x"0a400",-- 2624
x"0bb00",-- 2992
x"0b100",-- 2832
x"0a800",-- 2688
x"0c500",-- 3152
x"0e100",-- 3600
x"0e800",-- 3712
x"0f100",-- 3856
x"0f100",-- 3856
x"0f600",-- 3936
x"10500",-- 4176
x"10c00",-- 4288
x"11800",-- 4480
x"10e00",-- 4320
x"10f00",-- 4336
x"10700",-- 4208
x"0fd00",-- 4048
x"0b300",-- 2864
x"09500",-- 2384
x"0f400",-- 3904
x"10200",-- 4128
x"0c600",-- 3168
x"05700",-- 1392
x"01d00",-- 464
x"03800",-- 896
x"03a00",-- 928
x"04300",-- 1072
x"00500",-- 80
x"f7500",-- -2224
x"f2300",-- -3536
x"f3500",-- -3248
x"f7700",-- -2192
x"f5e00",-- -2592
x"ef200",-- -4320
x"ebf00",-- -5136
x"ea400",-- -5568
x"e9f00",-- -5648
x"ed200",-- -4832
x"efd00",-- -4144
x"ee200",-- -4576
x"ead00",-- -5424
x"ecd00",-- -4912
x"f0000",-- -4096
x"f0b00",-- -3920
x"f2400",-- -3520
x"f5b00",-- -2640
x"f7500",-- -2224
x"f6d00",-- -2352
x"f7500",-- -2224
x"f9e00",-- -1568
x"fc000",-- -1024
x"fe000",-- -512
x"01400",-- 320
x"02400",-- 576
x"00300",-- 48
x"fed00",-- -304
x"02600",-- 608
x"05a00",-- 1440
x"06200",-- 1568
x"05900",-- 1424
x"03a00",-- 928
x"01300",-- 304
x"01f00",-- 496
x"05b00",-- 1456
x"07100",-- 1808
x"04e00",-- 1248
x"00e00",-- 224
x"00900",-- 144
x"01300",-- 304
x"01800",-- 384
x"01d00",-- 464
x"00200",-- 32
x"fe000",-- -512
x"fbc00",-- -1088
x"fcb00",-- -848
x"fbc00",-- -1088
x"fb100",-- -1264
x"fa800",-- -1408
x"fb400",-- -1216
x"fb500",-- -1200
x"f8b00",-- -1872
x"f8700",-- -1936
x"f9700",-- -1680
x"faf00",-- -1296
x"fc600",-- -928
x"fcd00",-- -816
x"fbe00",-- -1056
x"fac00",-- -1344
x"fc000",-- -1024
x"00000",-- 0
x"01c00",-- 448
x"02200",-- 544
x"01500",-- 336
x"02300",-- 560
x"03c00",-- 960
x"05c00",-- 1472
x"08600",-- 2144
x"09000",-- 2304
x"08800",-- 2176
x"08b00",-- 2224
x"0a800",-- 2688
x"0b100",-- 2832
x"0bb00",-- 2992
x"0c400",-- 3136
x"0c900",-- 3216
x"0ce00",-- 3296
x"0b900",-- 2960
x"0ac00",-- 2752
x"0cc00",-- 3264
x"0d400",-- 3392
x"0d000",-- 3328
x"0cf00",-- 3312
x"0c300",-- 3120
x"0b600",-- 2912
x"0c300",-- 3120
x"0cb00",-- 3248
x"0bc00",-- 3008
x"08c00",-- 2240
x"05800",-- 1408
x"08300",-- 2096
x"0a500",-- 2640
x"0a200",-- 2592
x"06600",-- 1632
x"02200",-- 544
x"01100",-- 272
x"00700",-- 112
x"00d00",-- 208
x"00800",-- 128
x"fc300",-- -976
x"f6d00",-- -2352
x"f5200",-- -2784
x"f5900",-- -2672
x"f6100",-- -2544
x"f3000",-- -3328
x"f1600",-- -3744
x"f0800",-- -3968
x"eeb00",-- -4432
x"ef100",-- -4336
x"f0e00",-- -3872
x"f1700",-- -3728
x"f0900",-- -3952
x"f1f00",-- -3600
x"f3f00",-- -3088
x"f4c00",-- -2880
x"f4000",-- -3072
x"f5e00",-- -2592
x"f8200",-- -2016
x"f9b00",-- -1616
x"fac00",-- -1344
x"fc100",-- -1008
x"fc700",-- -912
x"fc300",-- -976
x"fe000",-- -512
x"00a00",-- 160
x"01800",-- 384
x"00700",-- 112
x"00400",-- 64
x"00900",-- 144
x"00d00",-- 208
x"00d00",-- 208
x"01a00",-- 416
x"00d00",-- 208
x"00600",-- 96
x"00700",-- 112
x"00300",-- 48
x"00400",-- 64
x"ff700",-- -144
x"ff200",-- -224
x"ff400",-- -192
x"ff500",-- -176
x"fdf00",-- -528
x"fdb00",-- -592
x"fdd00",-- -560
x"fcf00",-- -784
x"fd500",-- -688
x"fdb00",-- -592
x"fd700",-- -656
x"fd200",-- -736
x"fcd00",-- -816
x"fd800",-- -640
x"fe900",-- -368
x"fe200",-- -480
x"ff800",-- -128
x"ffd00",-- -48
x"00200",-- 32
x"00f00",-- 240
x"01900",-- 400
x"01600",-- 352
x"02900",-- 656
x"03f00",-- 1008
x"04000",-- 1024
x"05300",-- 1328
x"04400",-- 1088
x"04100",-- 1040
x"06900",-- 1680
x"04400",-- 1088
x"05800",-- 1408
x"08700",-- 2160
x"03e00",-- 992
x"05f00",-- 1520
x"06400",-- 1600
x"03900",-- 912
x"04800",-- 1152
x"04c00",-- 1216
x"05300",-- 1328
x"03e00",-- 992
x"02300",-- 560
x"03000",-- 768
x"03300",-- 816
x"03100",-- 784
x"01800",-- 384
x"02e00",-- 736
x"03500",-- 848
x"01a00",-- 416
x"02b00",-- 688
x"02a00",-- 672
x"01e00",-- 480
x"03900",-- 912
x"04200",-- 1056
x"02d00",-- 720
x"03a00",-- 928
x"03a00",-- 928
x"03300",-- 816
x"03f00",-- 1008
x"04500",-- 1104
x"05000",-- 1280
x"05600",-- 1376
x"04500",-- 1104
x"03b00",-- 944
x"03800",-- 896
x"02b00",-- 688
x"02800",-- 640
x"02400",-- 576
x"00f00",-- 240
x"00400",-- 64
x"ff800",-- -128
x"fe900",-- -368
x"fdd00",-- -560
x"fd300",-- -720
x"fc600",-- -928
x"fc000",-- -1024
x"fbd00",-- -1072
x"fb800",-- -1152
x"fb600",-- -1184
x"fb100",-- -1264
x"fab00",-- -1360
x"fac00",-- -1344
x"fb600",-- -1184
x"fb400",-- -1216
x"fbb00",-- -1104
x"fba00",-- -1120
x"fb600",-- -1184
x"fbb00",-- -1104
x"fb600",-- -1184
x"fb600",-- -1184
x"fb800",-- -1152
x"fb600",-- -1184
x"fb000",-- -1280
x"fb300",-- -1232
x"fac00",-- -1344
x"fa300",-- -1488
x"fad00",-- -1328
x"fa200",-- -1504
x"f9200",-- -1760
x"faf00",-- -1296
x"faf00",-- -1296
x"f9600",-- -1696
x"fac00",-- -1344
x"faf00",-- -1296
x"fa500",-- -1456
x"fb300",-- -1232
x"fb900",-- -1136
x"fbd00",-- -1072
x"fc800",-- -896
x"fd300",-- -720
x"fd600",-- -672
x"fdd00",-- -560
x"fe200",-- -480
x"feb00",-- -336
x"ff500",-- -176
x"ffd00",-- -48
x"00300",-- 48
x"00200",-- 32
x"00a00",-- 160
x"01000",-- 256
x"01600",-- 352
x"01c00",-- 448
x"01f00",-- 496
x"02100",-- 528
x"02400",-- 576
x"03100",-- 784
x"03700",-- 880
x"03700",-- 880
x"04000",-- 1024
x"04000",-- 1024
x"04100",-- 1040
x"04800",-- 1152
x"04700",-- 1136
x"04600",-- 1120
x"04800",-- 1152
x"04700",-- 1136
x"04700",-- 1136
x"04600",-- 1120
x"04300",-- 1072
x"03e00",-- 992
x"03900",-- 912
x"03700",-- 880
x"03400",-- 832
x"02f00",-- 752
x"02800",-- 640
x"02300",-- 560
x"01e00",-- 480
x"01800",-- 384
x"01700",-- 368
x"01200",-- 288
x"00f00",-- 240
x"00d00",-- 208
x"00800",-- 128
x"00700",-- 112
x"00300",-- 48
x"00100",-- 16
x"00600",-- 96
x"00200",-- 32
x"00000",-- 0
x"00500",-- 80
x"00200",-- 32
x"00500",-- 80
x"00800",-- 128
x"00c00",-- 192
x"01200",-- 288
x"01800",-- 384
x"01700",-- 368
x"02000",-- 512
x"02700",-- 624
x"02d00",-- 720
x"03a00",-- 928
x"03d00",-- 976
x"04200",-- 1056
x"04300",-- 1072
x"04100",-- 1040
x"04000",-- 1024
x"04000",-- 1024
x"03f00",-- 1008
x"03500",-- 848
x"03200",-- 800
x"02600",-- 608
x"01a00",-- 416
x"01400",-- 320
x"00500",-- 80
x"ffa00",-- -96
x"ff600",-- -160
x"fe400",-- -448
x"fe000",-- -512
x"fdc00",-- -576
x"fce00",-- -800
x"fd000",-- -768
x"fc800",-- -896
x"fc500",-- -944
x"fc200",-- -992
x"fbf00",-- -1040
x"fbc00",-- -1088
x"fbb00",-- -1104
x"fbb00",-- -1104
x"fb800",-- -1152
x"fba00",-- -1120
x"fb800",-- -1152
x"fb700",-- -1168
x"fb600",-- -1184
x"fb600",-- -1184
x"fb400",-- -1216
x"fb700",-- -1168
x"fb600",-- -1184
x"fb600",-- -1184
x"fbc00",-- -1088
x"fb900",-- -1136
x"fbb00",-- -1104
x"fbe00",-- -1056
x"fc000",-- -1024
x"fc600",-- -928
x"fca00",-- -864
x"fcf00",-- -784
x"fd200",-- -736
x"fd300",-- -720
x"fd900",-- -624
x"fe000",-- -512
x"fe900",-- -368
x"fec00",-- -320
x"ff000",-- -256
x"ff500",-- -176
x"ffa00",-- -96
x"00000",-- 0
x"00700",-- 112
x"00d00",-- 208
x"00d00",-- 208
x"01500",-- 336
x"01a00",-- 416
x"02000",-- 512
x"02400",-- 576
x"02600",-- 608
x"02b00",-- 688
x"03000",-- 768
x"03400",-- 832
x"03600",-- 864
x"03900",-- 912
x"03800",-- 896
x"03a00",-- 928
x"03d00",-- 976
x"03c00",-- 960
x"03900",-- 912
x"03700",-- 880
x"03500",-- 848
x"03400",-- 832
x"03200",-- 800
x"02e00",-- 736
x"02c00",-- 704
x"02600",-- 608
x"02200",-- 544
x"02200",-- 544
x"01f00",-- 496
x"01900",-- 400
x"01600",-- 352
x"01400",-- 320
x"01000",-- 256
x"00e00",-- 224
x"00d00",-- 208
x"00900",-- 144
x"00800",-- 128
x"00400",-- 64
x"00200",-- 32
x"00200",-- 32
x"00000",-- 0
x"fff00",-- -16
x"ffc00",-- -64
x"ffc00",-- -64
x"ffa00",-- -96
x"ff800",-- -128
x"ff800",-- -128
x"ff800",-- -128
x"ff600",-- -160
x"ff600",-- -160
x"ff500",-- -176
x"ff400",-- -192
x"ff400",-- -192
x"ff400",-- -192
x"ff400",-- -192
x"ff400",-- -192
x"ff500",-- -176
x"ff500",-- -176
x"ff600",-- -160
x"ff700",-- -144
x"ff800",-- -128
x"ff900",-- -112
x"ffd00",-- -48
x"ffe00",-- -32
x"00000",-- 0
x"00300",-- 48
x"00400",-- 64
x"00500",-- 80
x"00900",-- 144
x"00900",-- 144
x"00b00",-- 176
x"00b00",-- 176
x"00b00",-- 176
x"00b00",-- 176
x"00900",-- 144
x"00b00",-- 176
x"00700",-- 112
x"00700",-- 112
x"00400",-- 64
x"00100",-- 16
x"00200",-- 32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffb00",-- -80
x"ff900",-- -112
x"ff800",-- -128
x"ff500",-- -176
x"ff500",-- -176
x"ff200",-- -224
x"ff300",-- -208
x"ff100",-- -240
x"ff100",-- -240
x"ff000",-- -256
x"fee00",-- -288
x"fed00",-- -304
x"fec00",-- -320
x"fec00",-- -320
x"fea00",-- -352
x"fea00",-- -352
x"fe700",-- -400
x"fe500",-- -432
x"fe600",-- -416
x"fe500",-- -432
x"fe400",-- -448
x"fe400",-- -448
x"fe500",-- -432
x"fe500",-- -432
x"fe500",-- -432
x"fe700",-- -400
x"fe700",-- -400
x"fea00",-- -352
x"fec00",-- -320
x"fef00",-- -272
x"ff100",-- -240
x"ff300",-- -208
x"ff700",-- -144
x"ffa00",-- -96
x"ffe00",-- -32
x"00100",-- 16
x"00300",-- 48
x"00500",-- 80
x"00900",-- 144
x"00d00",-- 208
x"00f00",-- 240
x"01100",-- 272
x"01200",-- 288
x"01400",-- 320
x"01700",-- 368
x"01700",-- 368
x"01900",-- 400
x"01a00",-- 416
x"01a00",-- 416
x"01b00",-- 432
x"01c00",-- 448
x"01b00",-- 432
x"01b00",-- 432
x"01b00",-- 432
x"01a00",-- 416
x"01900",-- 400
x"01a00",-- 416
x"01a00",-- 416
x"01900",-- 400
x"01800",-- 384
x"01600",-- 352
x"01600",-- 352
x"01500",-- 336
x"01300",-- 304
x"01300",-- 304
x"01200",-- 288
x"00f00",-- 240
x"00c00",-- 192
x"00a00",-- 160
x"00900",-- 144
x"00600",-- 96
x"00400",-- 64
x"00200",-- 32
x"ffe00",-- -32
x"ffb00",-- -80
x"ff800",-- -128
x"ff700",-- -144
x"ff400",-- -192
x"ff300",-- -208
x"ff000",-- -256
x"fee00",-- -288
x"fec00",-- -320
x"feb00",-- -336
x"feb00",-- -336
x"fea00",-- -352
x"fe800",-- -384
x"fe800",-- -384
x"fe800",-- -384
x"fe800",-- -384
x"fe800",-- -384
x"fe900",-- -368
x"fea00",-- -352
x"fe900",-- -368
x"feb00",-- -336
x"fed00",-- -304
x"fee00",-- -288
x"fef00",-- -272
x"ff000",-- -256
x"ff200",-- -224
x"ff300",-- -208
x"ff400",-- -192
x"ff700",-- -144
x"ff800",-- -128
x"ff900",-- -112
x"ffa00",-- -96
x"ffb00",-- -80
x"ffd00",-- -48
x"fff00",-- -16
x"00000",-- 0
x"00200",-- 32
x"00200",-- 32
x"00300",-- 48
x"00500",-- 80
x"00600",-- 96
x"00700",-- 112
x"00700",-- 112
x"00800",-- 128
x"00900",-- 144
x"00900",-- 144
x"00a00",-- 160
x"00a00",-- 160
x"00b00",-- 176
x"00b00",-- 176
x"00b00",-- 176
x"00b00",-- 176
x"00a00",-- 160
x"00900",-- 144
x"00a00",-- 160
x"00900",-- 144
x"00800",-- 128
x"00800",-- 128
x"00600",-- 96
x"00500",-- 80
x"00500",-- 80
x"00500",-- 80
x"00300",-- 48
x"00300",-- 48
x"00300",-- 48
x"00200",-- 32
x"00300",-- 48
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"fff00",-- -16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffc00",-- -64
x"ffd00",-- -48
x"ffc00",-- -64
x"ffc00",-- -64
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffc00",-- -64
x"ffa00",-- -96
x"ffb00",-- -80
x"ffc00",-- -64
x"ffa00",-- -96
x"ffa00",-- -96
x"ff900",-- -112
x"ff800",-- -128
x"ff900",-- -112
x"ff900",-- -112
x"ff800",-- -128
x"ff800",-- -128
x"ff700",-- -144
x"ff700",-- -144
x"ff800",-- -128
x"ff800",-- -128
x"ff800",-- -128
x"ff800",-- -128
x"ff800",-- -128
x"ff800",-- -128
x"ff800",-- -128
x"ff800",-- -128
x"ff700",-- -144
x"ff700",-- -144
x"ff800",-- -128
x"ff800",-- -128
x"ff800",-- -128
x"ff800",-- -128
x"ff800",-- -128
x"ffa00",-- -96
x"ffa00",-- -96
x"ffb00",-- -80
x"ffb00",-- -80
x"ffb00",-- -80
x"ffc00",-- -64
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00300",-- 48
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00500",-- 80
x"00500",-- 80
x"00500",-- 80
x"00500",-- 80
x"00500",-- 80
x"00600",-- 96
x"00600",-- 96
x"00600",-- 96
x"00600",-- 96
x"00600",-- 96
x"00500",-- 80
x"00600",-- 96
x"00500",-- 80
x"00500",-- 80
x"00500",-- 80
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00300",-- 48
x"00300",-- 48
x"00300",-- 48
x"00300",-- 48
x"00300",-- 48
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"fff00",-- -16
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"ffc00",-- -64
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"ffd00",-- -48
x"ffe00",-- -32
x"ffc00",-- -64
x"ffe00",-- -32
x"ffa00",-- -96
x"ffb00",-- -80
x"ff200",-- -224
x"ff300",-- -208
x"fc300",-- -976
x"f8d00",-- -1840
x"00300",-- 48
x"04c00",-- 1216
x"00e00",-- 224
x"00400",-- 64
x"00500",-- 80
x"ff800",-- -128
x"01500",-- 336
x"01300",-- 304
x"00300",-- 48
x"ffa00",-- -96
x"00000",-- 0
x"00f00",-- 240
x"00800",-- 128
x"01400",-- 320
x"02300",-- 560
x"01800",-- 384
x"01400",-- 320
x"01200",-- 288
x"00000",-- 0
x"ffd00",-- -48
x"00200",-- 32
x"00300",-- 48
x"ffb00",-- -80
x"ffb00",-- -80
x"ff500",-- -176
x"ff700",-- -144
x"00600",-- 96
x"ff800",-- -128
x"ff700",-- -144
x"ffe00",-- -32
x"fff00",-- -16
x"ffc00",-- -64
x"01000",-- 256
x"01200",-- 288
x"ff800",-- -128
x"00600",-- 96
x"00300",-- 48
x"ff900",-- -112
x"02100",-- 528
x"00700",-- 112
x"ffc00",-- -64
x"01800",-- 384
x"ffe00",-- -32
x"01000",-- 256
x"fd200",-- -736
x"f7500",-- -2224
x"fff00",-- -16
x"03c00",-- 960
x"f9a00",-- -1632
x"fa300",-- -1488
x"02600",-- 608
x"01b00",-- 432
x"ff700",-- -144
x"ff700",-- -144
x"fed00",-- -304
x"ffd00",-- -48
x"02900",-- 656
x"00300",-- 48
x"fd900",-- -624
x"00800",-- 128
x"02c00",-- 704
x"01600",-- 352
x"01a00",-- 416
x"01b00",-- 432
x"01d00",-- 464
x"04400",-- 1088
x"01100",-- 272
x"00200",-- 32
x"04000",-- 1024
x"ffb00",-- -80
x"fe800",-- -384
x"02300",-- 560
x"ffd00",-- -48
x"fdc00",-- -576
x"01a00",-- 416
x"fed00",-- -304
x"fef00",-- -272
x"fff00",-- -16
x"ff300",-- -208
x"00e00",-- 224
x"fed00",-- -304
x"fed00",-- -304
x"00f00",-- 240
x"ffc00",-- -64
x"fed00",-- -304
x"fe800",-- -384
x"fe900",-- -368
x"fbf00",-- -1040
x"fb900",-- -1136
x"00200",-- 32
x"ff200",-- -224
x"ffa00",-- -96
x"fdd00",-- -560
x"fe700",-- -400
x"ff900",-- -112
x"00b00",-- 176
x"03a00",-- 928
x"01000",-- 256
x"fee00",-- -288
x"02300",-- 560
x"02c00",-- 704
x"ffb00",-- -80
x"00400",-- 64
x"04500",-- 1104
x"01a00",-- 416
x"01f00",-- 496
x"03100",-- 784
x"01900",-- 400
x"00900",-- 144
x"00a00",-- 160
x"02a00",-- 672
x"ff500",-- -176
x"ff800",-- -128
x"00c00",-- 192
x"fd200",-- -736
x"ff300",-- -208
x"ffd00",-- -48
x"fe200",-- -480
x"feb00",-- -336
x"fd000",-- -768
x"ff400",-- -192
x"00800",-- 128
x"ff100",-- -240
x"ff900",-- -112
x"fc700",-- -912
x"00b00",-- 176
x"fef00",-- -272
x"fe600",-- -416
x"01600",-- 352
x"fbb00",-- -1104
x"01700",-- 368
x"00700",-- 112
x"fea00",-- -352
x"03700",-- 880
x"ff900",-- -112
x"01c00",-- 448
x"03800",-- 896
x"fed00",-- -304
x"03300",-- 816
x"00600",-- 96
x"ff700",-- -144
x"01a00",-- 416
x"ff700",-- -144
x"03400",-- 832
x"ff800",-- -128
x"01a00",-- 416
x"02400",-- 576
x"00100",-- 16
x"00100",-- 16
x"02000",-- 512
x"fee00",-- -288
x"fef00",-- -272
x"03200",-- 800
x"fc700",-- -912
x"01f00",-- 496
x"fe000",-- -512
x"00e00",-- 224
x"ff900",-- -112
x"00800",-- 128
x"01000",-- 256
x"ff800",-- -128
x"00600",-- 96
x"ff800",-- -128
x"00900",-- 144
x"fd400",-- -704
x"03a00",-- 928
x"fd400",-- -704
x"fe700",-- -400
x"02500",-- 592
x"fc400",-- -960
x"fe000",-- -512
x"fd100",-- -752
x"fdf00",-- -528
x"02800",-- 640
x"fe900",-- -368
x"fee00",-- -288
x"04c00",-- 1216
x"fce00",-- -800
x"00e00",-- 224
x"01000",-- 256
x"fd100",-- -752
x"01500",-- 336
x"fe500",-- -432
x"02900",-- 656
x"00800",-- 128
x"faf00",-- -1296
x"05200",-- 1312
x"01b00",-- 432
x"fc300",-- -976
x"04400",-- 1088
x"02100",-- 528
x"fd700",-- -656
x"00800",-- 128
x"01500",-- 336
x"fbe00",-- -1056
x"05100",-- 1296
x"fdd00",-- -560
x"fdd00",-- -560
x"03e00",-- 992
x"fea00",-- -352
x"fe100",-- -496
x"fed00",-- -304
x"02d00",-- 720
x"fce00",-- -800
x"ff800",-- -128
x"03300",-- 816
x"fe400",-- -448
x"00f00",-- 240
x"01100",-- 272
x"fc400",-- -960
x"02d00",-- 720
x"fe900",-- -368
x"fd600",-- -672
x"04300",-- 1072
x"fe200",-- -480
x"ff200",-- -224
x"02900",-- 656
x"fbc00",-- -1088
x"01000",-- 256
x"04100",-- 1040
x"fb400",-- -1216
x"03500",-- 848
x"02400",-- 576
x"fba00",-- -1120
x"01c00",-- 448
x"00200",-- 32
x"fed00",-- -304
x"fef00",-- -272
x"01600",-- 352
x"00800",-- 128
x"fe900",-- -368
x"00400",-- 64
x"ff400",-- -192
x"fd600",-- -672
x"ff500",-- -176
x"fcc00",-- -832
x"00700",-- 112
x"00700",-- 112
x"fcc00",-- -832
x"fdb00",-- -592
x"01000",-- 256
x"fe400",-- -448
x"01f00",-- 496
x"00a00",-- 160
x"fe700",-- -400
x"03100",-- 784
x"ff800",-- -128
x"01f00",-- 496
x"01800",-- 384
x"ffd00",-- -48
x"01700",-- 368
x"03900",-- 912
x"02c00",-- 704
x"fe100",-- -496
x"02800",-- 640
x"fee00",-- -288
x"01a00",-- 416
x"00f00",-- 240
x"01500",-- 336
x"00d00",-- 208
x"fbe00",-- -1056
x"01800",-- 384
x"fff00",-- -16
x"fdf00",-- -528
x"ff600",-- -160
x"00600",-- 96
x"fb700",-- -1168
x"00000",-- 0
x"03200",-- 800
x"fc800",-- -896
x"fef00",-- -272
x"01600",-- 352
x"feb00",-- -336
x"00500",-- 80
x"03b00",-- 944
x"fd100",-- -752
x"fe100",-- -496
x"03d00",-- 976
x"fe900",-- -368
x"ffc00",-- -64
x"02800",-- 640
x"fef00",-- -272
x"fee00",-- -288
x"02d00",-- 720
x"ffc00",-- -64
x"00800",-- 128
x"01800",-- 384
x"fe200",-- -480
x"01800",-- 384
x"ffe00",-- -32
x"01100",-- 272
x"00b00",-- 176
x"fe500",-- -432
x"00e00",-- 224
x"00b00",-- 176
x"ffe00",-- -32
x"fbf00",-- -1040
x"03800",-- 896
x"ff300",-- -208
x"fad00",-- -1328
x"06400",-- 1600
x"fe000",-- -512
x"fc000",-- -1024
x"04200",-- 1056
x"fcc00",-- -832
x"ff900",-- -112
x"02e00",-- 736
x"ff900",-- -112
x"fe500",-- -432
x"00300",-- 48
x"01200",-- 288
x"fec00",-- -320
x"00200",-- 32
x"ff900",-- -112
x"01d00",-- 464
x"fe400",-- -448
x"ff900",-- -112
x"02f00",-- 752
x"fd200",-- -736
x"ffd00",-- -48
x"02c00",-- 704
x"ff200",-- -224
x"fda00",-- -608
x"04200",-- 1056
x"00400",-- 64
x"fc300",-- -976
x"00f00",-- 240
x"01d00",-- 464
x"fec00",-- -320
x"ff500",-- -176
x"02300",-- 560
x"fea00",-- -352
x"00c00",-- 192
x"00a00",-- 160
x"fe300",-- -464
x"01c00",-- 448
x"00900",-- 144
x"fdc00",-- -576
x"01800",-- 384
x"00100",-- 16
x"ff600",-- -160
x"00a00",-- 160
x"fff00",-- -16
x"fe100",-- -496
x"03200",-- 800
x"ff800",-- -128
x"fcb00",-- -848
x"03b00",-- 944
x"fc600",-- -928
x"fed00",-- -304
x"04000",-- 1024
x"fc000",-- -1024
x"fd900",-- -624
x"04800",-- 1152
x"fd500",-- -688
x"fe700",-- -400
x"00700",-- 112
x"01100",-- 272
x"00a00",-- 160
x"fdd00",-- -560
x"00000",-- 0
x"01d00",-- 464
x"fed00",-- -304
x"fed00",-- -304
x"02400",-- 576
x"ff500",-- -176
x"00100",-- 16
x"02b00",-- 688
x"fee00",-- -288
x"fea00",-- -352
x"04700",-- 1136
x"fc000",-- -1024
x"ffd00",-- -48
x"03300",-- 816
x"fd400",-- -704
x"00600",-- 96
x"00200",-- 32
x"ff300",-- -208
x"fd800",-- -640
x"02400",-- 576
x"00b00",-- 176
x"fb200",-- -1248
x"06200",-- 1568
x"fe900",-- -368
x"fb400",-- -1216
x"05900",-- 1424
x"fcd00",-- -816
x"ff400",-- -192
x"02000",-- 512
x"fea00",-- -352
x"02200",-- 544
x"fc300",-- -976
x"00f00",-- 240
x"03900",-- 912
x"fb900",-- -1136
x"01c00",-- 448
x"02300",-- 560
x"fed00",-- -304
x"01500",-- 336
x"ffd00",-- -48
x"fe000",-- -512
x"01f00",-- 496
x"00100",-- 16
x"fd200",-- -736
x"03100",-- 784
x"fe100",-- -496
x"fd900",-- -624
x"02000",-- 512
x"00900",-- 144
x"ffc00",-- -64
x"ff500",-- -176
x"00200",-- 32
x"00c00",-- 192
x"00100",-- 16
x"fc700",-- -912
x"02500",-- 592
x"02700",-- 624
x"fa600",-- -1440
x"02800",-- 640
x"04d00",-- 1232
x"fa200",-- -1504
x"00900",-- 144
x"03800",-- 896
x"fd000",-- -768
x"01c00",-- 448
x"00400",-- 64
x"fb800",-- -1152
x"01a00",-- 416
x"03c00",-- 960
x"fb400",-- -1216
x"01e00",-- 480
x"03600",-- 864
x"faa00",-- -1376
x"03000",-- 768
x"00800",-- 128
x"fe400",-- -448
x"01700",-- 368
x"fe800",-- -384
x"fe200",-- -480
x"02400",-- 576
x"04200",-- 1056
x"fbe00",-- -1056
x"fed00",-- -304
x"03800",-- 896
x"fdc00",-- -576
x"00500",-- 80
x"03a00",-- 928
x"fbc00",-- -1088
x"01b00",-- 432
x"01800",-- 384
x"fef00",-- -272
x"02700",-- 624
x"fcb00",-- -848
x"00100",-- 16
x"02a00",-- 672
x"fe800",-- -384
x"02900",-- 656
x"feb00",-- -336
x"ff100",-- -240
x"00f00",-- 240
x"fec00",-- -320
x"03300",-- 816
x"ff400",-- -192
x"fee00",-- -288
x"fe000",-- -512
x"01600",-- 352
x"00100",-- 16
x"fc700",-- -912
x"00200",-- 32
x"02100",-- 528
x"fe100",-- -496
x"fac00",-- -1344
x"03d00",-- 976
x"fe100",-- -496
x"ffd00",-- -48
x"fe700",-- -400
x"ff800",-- -128
x"05800",-- 1408
x"fcb00",-- -848
x"01200",-- 288
x"ff200",-- -224
x"00100",-- 16
x"03b00",-- 944
x"fe800",-- -384
x"02500",-- 592
x"02400",-- 576
x"fe400",-- -448
x"03a00",-- 928
x"fdd00",-- -560
x"01400",-- 320
x"04c00",-- 1216
x"fcb00",-- -848
x"ffc00",-- -64
x"04e00",-- 1248
x"ff800",-- -128
x"fc700",-- -912
x"01500",-- 336
x"ff500",-- -176
x"00500",-- 80
x"01700",-- 368
x"fdd00",-- -560
x"01300",-- 304
x"02300",-- 560
x"fc400",-- -960
x"01e00",-- 480
x"02400",-- 576
x"fef00",-- -272
x"00000",-- 0
x"01800",-- 384
x"01a00",-- 416
x"fe400",-- -448
x"00200",-- 32
x"01f00",-- 496
x"02000",-- 512
x"fd500",-- -688
x"02c00",-- 704
x"02700",-- 624
x"fe300",-- -464
x"ff800",-- -128
x"00f00",-- 240
x"01d00",-- 464
x"fcf00",-- -784
x"02700",-- 624
x"03c00",-- 960
x"fe000",-- -512
x"fc200",-- -992
x"00b00",-- 176
x"03200",-- 800
x"fe500",-- -432
x"feb00",-- -336
x"01100",-- 272
x"ff900",-- -112
x"ffd00",-- -48
x"fe200",-- -480
x"01600",-- 352
x"02400",-- 576
x"fae00",-- -1312
x"ffc00",-- -64
x"05100",-- 1296
x"ff300",-- -208
x"fdd00",-- -560
x"01a00",-- 416
x"00000",-- 0
x"00300",-- 48
x"01a00",-- 416
x"01100",-- 272
x"01900",-- 400
x"fd800",-- -640
x"fe500",-- -432
x"05700",-- 1392
x"fed00",-- -304
x"fe400",-- -448
x"02300",-- 560
x"fd000",-- -768
x"01400",-- 320
x"00a00",-- 160
x"fda00",-- -608
x"01a00",-- 416
x"fe600",-- -416
x"ff100",-- -240
x"03600",-- 864
x"fec00",-- -320
x"fe700",-- -400
x"ff000",-- -256
x"01400",-- 320
x"01c00",-- 448
x"ffc00",-- -64
x"fe400",-- -448
x"ff400",-- -192
x"ff800",-- -128
x"ff700",-- -144
x"03700",-- 880
x"fe100",-- -496
x"ff800",-- -128
x"01900",-- 400
x"fb200",-- -1248
x"03c00",-- 960
x"02800",-- 640
x"fa200",-- -1504
x"04500",-- 1104
x"01300",-- 304
x"fbd00",-- -1072
x"01400",-- 320
x"01900",-- 400
x"fc200",-- -992
x"03b00",-- 944
x"01d00",-- 464
x"f8e00",-- -1824
x"02500",-- 592
x"05000",-- 1280
x"fd900",-- -624
x"fed00",-- -304
x"01000",-- 256
x"fe100",-- -496
x"02000",-- 512
x"ff700",-- -144
x"ff300",-- -208
x"02d00",-- 720
x"fb700",-- -1168
x"fdd00",-- -560
x"08c00",-- 2240
x"fc400",-- -960
x"f8400",-- -1984
x"06500",-- 1616
x"fea00",-- -352
x"fd400",-- -704
x"04500",-- 1104
x"fc700",-- -912
x"fca00",-- -864
x"03d00",-- 976
x"ff400",-- -192
x"03700",-- 880
x"00000",-- 0
x"f8200",-- -2016
x"03000",-- 768
x"03c00",-- 960
x"fee00",-- -288
x"fec00",-- -320
x"02400",-- 576
x"01800",-- 384
x"fb900",-- -1136
x"00000",-- 0
x"05600",-- 1376
x"ffc00",-- -64
x"fb900",-- -1136
x"01d00",-- 464
x"03800",-- 896
x"ffa00",-- -96
x"fc000",-- -1024
x"fe400",-- -448
x"03d00",-- 976
x"ff000",-- -256
x"fd200",-- -736
x"02900",-- 656
x"ff500",-- -176
x"fcc00",-- -832
x"00a00",-- 160
x"02c00",-- 704
x"00100",-- 16
x"fac00",-- -1344
x"01a00",-- 416
x"04500",-- 1104
x"fb900",-- -1136
x"fdd00",-- -560
x"04e00",-- 1248
x"00100",-- 16
x"fb300",-- -1232
x"01000",-- 256
x"04900",-- 1168
x"fdd00",-- -560
x"fb600",-- -1184
x"03600",-- 864
x"02e00",-- 736
x"fef00",-- -272
x"fdc00",-- -576
x"ff500",-- -176
x"03f00",-- 1008
x"fca00",-- -864
x"fd600",-- -672
x"04b00",-- 1200
x"00600",-- 96
x"f9c00",-- -1600
x"00400",-- 64
x"05400",-- 1344
x"ff100",-- -240
x"fde00",-- -544
x"fd900",-- -624
x"00f00",-- 240
x"02400",-- 576
x"fd000",-- -768
x"00f00",-- 240
x"05700",-- 1392
x"fac00",-- -1344
x"faa00",-- -1376
x"07800",-- 1920
x"03500",-- 848
x"f9700",-- -1680
x"02800",-- 640
x"02000",-- 512
x"fc000",-- -1024
x"00a00",-- 160
x"00200",-- 32
x"ffb00",-- -80
x"01900",-- 400
x"fff00",-- -16
x"fff00",-- -16
x"01a00",-- 416
x"fde00",-- -544
x"fdf00",-- -528
x"00e00",-- 224
x"02800",-- 640
x"fef00",-- -272
x"fd900",-- -624
x"02100",-- 528
x"01500",-- 336
x"fbf00",-- -1040
x"00b00",-- 176
x"05900",-- 1424
x"ff100",-- -240
x"fbc00",-- -1088
x"01f00",-- 496
x"02d00",-- 720
x"fb500",-- -1200
x"01400",-- 320
x"02e00",-- 736
x"fd600",-- -672
x"00200",-- 32
x"fe700",-- -400
x"01600",-- 352
x"03600",-- 864
x"fbc00",-- -1088
x"ffb00",-- -80
x"01d00",-- 464
x"fc700",-- -912
x"ff900",-- -112
x"02a00",-- 672
x"fef00",-- -272
x"fee00",-- -288
x"ffe00",-- -32
x"ff300",-- -208
x"03c00",-- 960
x"fe400",-- -448
x"fac00",-- -1344
x"05d00",-- 1488
x"02500",-- 592
x"fa800",-- -1408
x"02000",-- 512
x"02900",-- 656
x"fd100",-- -752
x"02400",-- 576
x"02400",-- 576
x"fe000",-- -512
x"00000",-- 0
x"fe100",-- -496
x"ff700",-- -144
x"04600",-- 1120
x"00d00",-- 208
x"ff300",-- -208
x"01200",-- 288
x"fde00",-- -544
x"00000",-- 0
x"01200",-- 288
x"fdc00",-- -576
x"ff800",-- -128
x"ffc00",-- -64
x"00700",-- 112
x"01200",-- 288
x"ffe00",-- -32
x"ff500",-- -176
x"fe200",-- -480
x"ffb00",-- -80
x"01800",-- 384
x"01600",-- 352
x"fe600",-- -416
x"00400",-- 64
x"00a00",-- 160
x"00400",-- 64
x"02d00",-- 720
x"ffb00",-- -80
x"fe900",-- -368
x"ff400",-- -192
x"02000",-- 512
x"00b00",-- 176
x"00400",-- 64
x"02100",-- 528
x"fcd00",-- -816
x"fe600",-- -416
x"03400",-- 832
x"01c00",-- 448
x"fe800",-- -384
x"ff900",-- -112
x"ff700",-- -144
x"fe800",-- -384
x"ff700",-- -144
x"ff400",-- -192
x"00900",-- 144
x"fef00",-- -272
x"01c00",-- 448
x"00500",-- 80
x"fc300",-- -976
x"00800",-- 128
x"ff300",-- -208
x"fde00",-- -544
x"03100",-- 784
x"02700",-- 624
x"fed00",-- -304
x"fe300",-- -464
x"ffc00",-- -64
x"01600",-- 352
x"fea00",-- -352
x"ffa00",-- -96
x"01d00",-- 464
x"00700",-- 112
x"ff300",-- -208
x"01900",-- 400
x"fe800",-- -384
x"fec00",-- -320
x"02400",-- 576
x"fe400",-- -448
x"00d00",-- 208
x"01600",-- 352
x"fee00",-- -288
x"00300",-- 48
x"fe000",-- -512
x"fff00",-- -16
x"ffe00",-- -32
x"fde00",-- -544
x"00500",-- 80
x"01400",-- 320
x"ffd00",-- -48
x"fd900",-- -624
x"ff200",-- -224
x"ffb00",-- -80
x"ff100",-- -240
x"ffa00",-- -96
x"fef00",-- -272
x"00200",-- 32
x"00300",-- 48
x"fef00",-- -272
x"fed00",-- -304
x"01000",-- 256
x"ff300",-- -208
x"fde00",-- -544
x"04100",-- 1040
x"02300",-- 560
x"fc700",-- -912
x"fe200",-- -480
x"00800",-- 128
x"00c00",-- 192
x"ff100",-- -240
x"ff800",-- -128
x"02900",-- 656
x"ffa00",-- -96
x"fcd00",-- -816
x"01f00",-- 496
x"01a00",-- 416
x"fe500",-- -432
x"fe700",-- -400
x"01000",-- 256
x"01800",-- 384
x"ff200",-- -224
x"01300",-- 304
x"fec00",-- -320
x"ffc00",-- -64
x"02a00",-- 672
x"fde00",-- -544
x"fee00",-- -288
x"02a00",-- 672
x"feb00",-- -336
x"ff900",-- -112
x"03300",-- 816
x"ff600",-- -160
x"fed00",-- -304
x"00300",-- 48
x"00d00",-- 208
x"ffa00",-- -96
x"ff600",-- -160
x"02300",-- 560
x"ff800",-- -128
x"fd400",-- -704
x"01e00",-- 480
x"01d00",-- 464
x"ffa00",-- -96
x"01400",-- 320
x"00100",-- 16
x"feb00",-- -336
x"01b00",-- 432
x"00500",-- 80
x"feb00",-- -336
x"01d00",-- 464
x"02e00",-- 736
x"ff900",-- -112
x"fec00",-- -320
x"04200",-- 1056
x"00400",-- 64
x"fe100",-- -496
x"03700",-- 880
x"02700",-- 624
x"fff00",-- -16
x"00500",-- 80
x"01e00",-- 480
x"00900",-- 144
x"ff400",-- -192
x"02b00",-- 688
x"03400",-- 832
x"ff100",-- -240
x"fef00",-- -272
x"02400",-- 576
x"01500",-- 336
x"feb00",-- -336
x"00500",-- 80
x"02200",-- 544
x"00200",-- 32
x"ff000",-- -256
x"01000",-- 256
x"00e00",-- 224
x"ff400",-- -192
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffa00",-- -96
x"00e00",-- 224
x"00900",-- 144
x"ffe00",-- -32
x"00200",-- 32
x"ff800",-- -128
x"fee00",-- -288
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"fe900",-- -368
x"fdd00",-- -560
x"ff800",-- -128
x"fed00",-- -304
x"fe100",-- -496
x"fe700",-- -400
x"ff900",-- -112
x"fe500",-- -432
x"fbe00",-- -1056
x"fe500",-- -432
x"fe800",-- -384
x"fcb00",-- -848
x"fdf00",-- -528
x"fea00",-- -352
x"fd400",-- -704
x"fbb00",-- -1104
x"fc900",-- -880
x"fed00",-- -304
x"fd400",-- -704
x"fc800",-- -896
x"fe500",-- -432
x"fed00",-- -304
x"fcd00",-- -816
x"fc800",-- -896
x"ff400",-- -192
x"ff000",-- -256
x"fc600",-- -928
x"fc500",-- -944
x"00000",-- 0
x"00900",-- 144
x"fba00",-- -1120
x"fd600",-- -672
x"01f00",-- 496
x"fef00",-- -272
x"fcc00",-- -832
x"ffa00",-- -96
x"02300",-- 560
x"ffd00",-- -48
x"fd500",-- -688
x"00300",-- 48
x"02e00",-- 736
x"ff000",-- -256
x"ff800",-- -128
x"02c00",-- 704
x"00e00",-- 224
x"ff300",-- -208
x"01000",-- 256
x"06600",-- 1632
x"02100",-- 528
x"fef00",-- -272
x"06400",-- 1600
x"06b00",-- 1712
x"fec00",-- -320
x"01b00",-- 432
x"09700",-- 2416
x"03e00",-- 992
x"00800",-- 128
x"06a00",-- 1696
x"07900",-- 1936
x"04400",-- 1088
x"03800",-- 896
x"04100",-- 1040
x"05500",-- 1360
x"05e00",-- 1504
x"05800",-- 1408
x"07f00",-- 2032
x"08300",-- 2096
x"03100",-- 784
x"02700",-- 624
x"06a00",-- 1696
x"06700",-- 1648
x"03d00",-- 976
x"04c00",-- 1216
x"08400",-- 2112
x"06000",-- 1536
x"01300",-- 304
x"05d00",-- 1488
x"08900",-- 2192
x"02f00",-- 752
x"01800",-- 384
x"06200",-- 1568
x"04800",-- 1152
x"00500",-- 80
x"01600",-- 352
x"02f00",-- 752
x"00c00",-- 192
x"fd400",-- -704
x"fdb00",-- -592
x"fef00",-- -272
x"fc800",-- -896
x"f9b00",-- -1616
x"fb700",-- -1168
x"fae00",-- -1312
x"f7000",-- -2304
x"f7b00",-- -2128
x"f9800",-- -1664
x"f7f00",-- -2064
x"f6200",-- -2528
x"f5e00",-- -2592
x"f6a00",-- -2400
x"f6d00",-- -2352
x"f5900",-- -2672
x"f6500",-- -2480
x"f7f00",-- -2064
x"f6800",-- -2432
x"f5f00",-- -2576
x"f8200",-- -2016
x"f9700",-- -1680
x"f8300",-- -2000
x"f7f00",-- -2064
x"f9b00",-- -1616
x"f9f00",-- -1552
x"f9900",-- -1648
x"fb500",-- -1200
x"fb800",-- -1152
x"fab00",-- -1360
x"fad00",-- -1328
x"fb800",-- -1152
x"fca00",-- -864
x"fc800",-- -896
x"fbd00",-- -1072
x"fc800",-- -896
x"fca00",-- -864
x"fd100",-- -752
x"fdb00",-- -592
x"fd600",-- -672
x"fd300",-- -720
x"fcf00",-- -784
x"ffa00",-- -96
x"fea00",-- -352
x"fd600",-- -672
x"00f00",-- 240
x"01300",-- 304
x"feb00",-- -336
x"01700",-- 368
x"02f00",-- 752
x"01500",-- 336
x"03a00",-- 928
x"03100",-- 784
x"04700",-- 1136
x"05f00",-- 1520
x"05700",-- 1392
x"07600",-- 1888
x"08600",-- 2144
x"07700",-- 1904
x"05b00",-- 1456
x"09000",-- 2304
x"0ba00",-- 2976
x"08600",-- 2144
x"07100",-- 1808
x"0cf00",-- 3312
x"0e500",-- 3664
x"06f00",-- 1776
x"07d00",-- 2000
x"0ee00",-- 3808
x"0a900",-- 2704
x"07b00",-- 1968
x"0c900",-- 3216
x"0d800",-- 3456
x"0b300",-- 2864
x"09d00",-- 2512
x"0b900",-- 2960
x"0ca00",-- 3232
x"0ab00",-- 2736
x"09000",-- 2304
x"09400",-- 2368
x"0a000",-- 2560
x"07700",-- 1904
x"04400",-- 1088
x"05900",-- 1424
x"04e00",-- 1248
x"00e00",-- 224
x"00900",-- 144
x"02000",-- 512
x"ff600",-- -160
x"faa00",-- -1376
x"f9c00",-- -1600
x"fa900",-- -1392
x"f7900",-- -2160
x"f4300",-- -3024
x"f5c00",-- -2624
x"f6400",-- -2496
x"f3000",-- -3328
x"f2000",-- -3584
x"f3b00",-- -3152
x"f3900",-- -3184
x"f1800",-- -3712
x"f3100",-- -3312
x"f6300",-- -2512
x"f6900",-- -2416
x"f5e00",-- -2592
x"f7900",-- -2160
x"f9f00",-- -1552
x"f9600",-- -1696
x"fa300",-- -1488
x"fce00",-- -800
x"fe000",-- -512
x"fd600",-- -672
x"fdb00",-- -592
x"fee00",-- -288
x"fed00",-- -304
x"fe500",-- -432
x"fe600",-- -416
x"ff000",-- -256
x"ff100",-- -240
x"fdc00",-- -576
x"fd700",-- -656
x"fd300",-- -720
x"fb500",-- -1200
x"fa800",-- -1408
x"fa400",-- -1472
x"fa200",-- -1504
x"f9f00",-- -1552
x"f9500",-- -1712
x"f8a00",-- -1888
x"f8400",-- -1984
x"f7f00",-- -2064
x"f8800",-- -1920
x"fa700",-- -1424
x"fb900",-- -1136
x"fb500",-- -1200
x"fc200",-- -992
x"fd300",-- -720
x"fd800",-- -640
x"ff800",-- -128
x"00b00",-- 176
x"01600",-- 352
x"02c00",-- 704
x"03200",-- 800
x"05f00",-- 1520
x"06300",-- 1584
x"02c00",-- 704
x"05500",-- 1360
x"0a100",-- 2576
x"05d00",-- 1488
x"05800",-- 1408
x"0b900",-- 2960
x"07d00",-- 2000
x"04400",-- 1088
x"08300",-- 2096
x"0a100",-- 2576
x"06900",-- 1680
x"05a00",-- 1440
x"08a00",-- 2208
x"08d00",-- 2256
x"06a00",-- 1696
x"03c00",-- 960
x"07100",-- 1808
x"0a600",-- 2656
x"07200",-- 1824
x"06200",-- 1568
x"0aa00",-- 2720
x"0ae00",-- 2784
x"07e00",-- 2016
x"08c00",-- 2240
x"0aa00",-- 2720
x"0c400",-- 3136
x"0ab00",-- 2736
x"0ae00",-- 2784
x"0d700",-- 3440
x"0b000",-- 2816
x"07700",-- 1904
x"07400",-- 1856
x"07c00",-- 1984
x"06400",-- 1600
x"04c00",-- 1216
x"05100",-- 1296
x"03600",-- 864
x"00400",-- 64
x"fe800",-- -384
x"fe200",-- -480
x"fb700",-- -1168
x"f7200",-- -2272
x"f6900",-- -2416
x"f7b00",-- -2128
x"f5600",-- -2720
x"f2b00",-- -3408
x"f2f00",-- -3344
x"f1d00",-- -3632
x"f0100",-- -4080
x"f0b00",-- -3920
x"f3600",-- -3232
x"f3e00",-- -3104
x"f3600",-- -3232
x"f4a00",-- -2912
x"f7100",-- -2288
x"f8000",-- -2048
x"f8000",-- -2048
x"fa300",-- -1488
x"fc200",-- -992
x"fcc00",-- -832
x"fde00",-- -544
x"ffe00",-- -32
x"00600",-- 96
x"ffe00",-- -32
x"00400",-- 64
x"00f00",-- 240
x"00f00",-- 240
x"00500",-- 80
x"00500",-- 80
x"00500",-- 80
x"ff300",-- -208
x"fd500",-- -688
x"fcb00",-- -848
x"fc300",-- -976
x"fac00",-- -1344
x"fa400",-- -1472
x"fa800",-- -1408
x"fa300",-- -1488
x"f8d00",-- -1840
x"f7f00",-- -2064
x"f8600",-- -1952
x"f8e00",-- -1824
x"f8300",-- -2000
x"f8100",-- -2032
x"f9900",-- -1648
x"fb200",-- -1248
x"fc500",-- -944
x"fd000",-- -768
x"fd700",-- -656
x"fe000",-- -512
x"ff600",-- -160
x"00f00",-- 240
x"02100",-- 528
x"02300",-- 560
x"02c00",-- 704
x"03d00",-- 976
x"04800",-- 1152
x"05500",-- 1360
x"05d00",-- 1488
x"05e00",-- 1504
x"04400",-- 1088
x"04500",-- 1104
x"08300",-- 2096
x"08900",-- 2192
x"02500",-- 592
x"04a00",-- 1184
x"0a400",-- 2624
x"05100",-- 1296
x"01d00",-- 464
x"07500",-- 1872
x"09a00",-- 2464
x"03c00",-- 960
x"02100",-- 528
x"09a00",-- 2464
x"09000",-- 2304
x"02900",-- 656
x"05900",-- 1424
x"0bd00",-- 3024
x"09200",-- 2336
x"05d00",-- 1488
x"0ab00",-- 2736
x"0bb00",-- 2992
x"09000",-- 2304
x"0a500",-- 2640
x"0b000",-- 2816
x"0a600",-- 2656
x"0a300",-- 2608
x"07f00",-- 2032
x"05e00",-- 1504
x"06d00",-- 1744
x"07000",-- 1792
x"05000",-- 1280
x"04800",-- 1152
x"04900",-- 1168
x"02000",-- 512
x"ff100",-- -240
x"ff400",-- -192
x"fe100",-- -496
x"f9e00",-- -1568
x"f8a00",-- -1888
x"fa400",-- -1472
x"f8300",-- -2000
x"f5200",-- -2784
x"f6200",-- -2528
x"f5c00",-- -2624
x"f2900",-- -3440
x"f2500",-- -3504
x"f5500",-- -2736
x"f5b00",-- -2640
x"f4b00",-- -2896
x"f5f00",-- -2576
x"f8300",-- -2000
x"f8400",-- -1984
x"f7900",-- -2160
x"f9d00",-- -1584
x"fb600",-- -1184
x"fb500",-- -1200
x"fc500",-- -944
x"ff100",-- -240
x"ffa00",-- -96
x"fed00",-- -304
x"ff800",-- -128
x"00600",-- 96
x"00300",-- 48
x"ff700",-- -144
x"00300",-- 48
x"00900",-- 144
x"ffb00",-- -80
x"fe800",-- -384
x"fdb00",-- -592
x"fcc00",-- -832
x"fb900",-- -1136
x"fc000",-- -1024
x"fc700",-- -912
x"fbf00",-- -1040
x"fac00",-- -1344
x"fa100",-- -1520
x"fa200",-- -1504
x"fa800",-- -1408
x"fa600",-- -1440
x"fad00",-- -1328
x"fc000",-- -1024
x"fc000",-- -1024
x"fc900",-- -880
x"fdc00",-- -576
x"fd500",-- -688
x"fd300",-- -720
x"fe700",-- -400
x"00300",-- 48
x"01d00",-- 464
x"02200",-- 544
x"01900",-- 400
x"01e00",-- 480
x"02d00",-- 720
x"02200",-- 544
x"02400",-- 576
x"02e00",-- 736
x"03400",-- 832
x"04700",-- 1136
x"03300",-- 816
x"02300",-- 560
x"03b00",-- 944
x"04300",-- 1072
x"01d00",-- 464
x"00f00",-- 240
x"04d00",-- 1232
x"05500",-- 1360
x"01500",-- 336
x"02900",-- 656
x"04c00",-- 1216
x"03800",-- 896
x"02700",-- 624
x"04100",-- 1040
x"05300",-- 1328
x"03900",-- 912
x"03e00",-- 992
x"05600",-- 1376
x"05100",-- 1296
x"04200",-- 1056
x"04a00",-- 1184
x"06600",-- 1632
x"05500",-- 1360
x"05500",-- 1360
x"07900",-- 1936
x"06700",-- 1648
x"05200",-- 1312
x"06d00",-- 1744
x"07800",-- 1920
x"05700",-- 1392
x"05000",-- 1280
x"05e00",-- 1504
x"06500",-- 1616
x"06400",-- 1600
x"06300",-- 1584
x"06400",-- 1600
x"05400",-- 1344
x"03e00",-- 992
x"03400",-- 832
x"02600",-- 608
x"01400",-- 320
x"00800",-- 128
x"ffc00",-- -64
x"fea00",-- -352
x"fdd00",-- -560
x"fd400",-- -704
x"fc400",-- -960
x"fb200",-- -1248
x"fa700",-- -1424
x"fa300",-- -1488
x"fa100",-- -1520
x"fa200",-- -1504
x"fa300",-- -1488
x"fa100",-- -1520
x"f9b00",-- -1616
x"f9900",-- -1648
x"fa200",-- -1504
x"fa800",-- -1408
x"fac00",-- -1344
x"fb800",-- -1152
x"fc000",-- -1024
x"fc000",-- -1024
x"fc700",-- -912
x"fca00",-- -864
x"fc400",-- -960
x"fbf00",-- -1040
x"fba00",-- -1120
x"fbf00",-- -1040
x"fbd00",-- -1072
x"fb900",-- -1136
x"fb900",-- -1136
x"fb800",-- -1152
x"fb500",-- -1200
x"fb500",-- -1200
x"fbf00",-- -1040
x"fbb00",-- -1104
x"fbd00",-- -1072
x"fc200",-- -992
x"fc500",-- -944
x"fca00",-- -864
x"fce00",-- -800
x"fcf00",-- -784
x"fcc00",-- -832
x"fdb00",-- -592
x"fec00",-- -320
x"ff500",-- -176
x"ff600",-- -160
x"ff100",-- -240
x"ff600",-- -160
x"ff900",-- -112
x"ffb00",-- -80
x"fff00",-- -16
x"00200",-- 32
x"ffd00",-- -48
x"ffd00",-- -48
x"00700",-- 112
x"00b00",-- 176
x"00900",-- 144
x"00400",-- 64
x"00d00",-- 208
x"01300",-- 304
x"01300",-- 304
x"01a00",-- 416
x"02400",-- 576
x"02300",-- 560
x"01f00",-- 496
x"02700",-- 624
x"02f00",-- 752
x"02b00",-- 688
x"02a00",-- 672
x"02f00",-- 752
x"03100",-- 784
x"02d00",-- 720
x"03100",-- 784
x"03200",-- 800
x"03000",-- 768
x"02e00",-- 736
x"02c00",-- 704
x"02c00",-- 704
x"02900",-- 656
x"02b00",-- 688
x"02700",-- 624
x"02600",-- 608
x"02800",-- 640
x"02600",-- 608
x"02700",-- 624
x"02900",-- 656
x"02c00",-- 704
x"02b00",-- 688
x"02f00",-- 752
x"03500",-- 848
x"03a00",-- 928
x"03e00",-- 992
x"04200",-- 1056
x"04a00",-- 1184
x"04c00",-- 1216
x"05200",-- 1312
x"05b00",-- 1456
x"05f00",-- 1520
x"05e00",-- 1504
x"05e00",-- 1504
x"05e00",-- 1504
x"05800",-- 1408
x"05000",-- 1280
x"04c00",-- 1216
x"04600",-- 1120
x"03a00",-- 928
x"03000",-- 768
x"02800",-- 640
x"01d00",-- 464
x"01000",-- 256
x"00200",-- 32
x"ff900",-- -112
x"fed00",-- -304
x"fe500",-- -432
x"fdf00",-- -528
x"fda00",-- -608
x"fd400",-- -704
x"fcb00",-- -848
x"fc900",-- -880
x"fc500",-- -944
x"fbc00",-- -1088
x"fb600",-- -1184
x"fb500",-- -1200
x"faf00",-- -1296
x"fac00",-- -1344
x"fa800",-- -1408
x"fa800",-- -1408
x"fa300",-- -1488
x"f9c00",-- -1600
x"f9900",-- -1648
x"f9900",-- -1648
x"f9800",-- -1664
x"f9400",-- -1728
x"f9600",-- -1696
x"f9b00",-- -1616
x"f9a00",-- -1632
x"f9a00",-- -1632
x"f9e00",-- -1568
x"fa300",-- -1488
x"fa700",-- -1424
x"faa00",-- -1376
x"fb400",-- -1216
x"fbb00",-- -1104
x"fbf00",-- -1040
x"fc600",-- -928
x"fd100",-- -752
x"fd600",-- -672
x"fdc00",-- -576
x"fe500",-- -432
x"fea00",-- -352
x"fef00",-- -272
x"ff500",-- -176
x"ffb00",-- -80
x"fff00",-- -16
x"00200",-- 32
x"00600",-- 96
x"00900",-- 144
x"00f00",-- 240
x"01300",-- 304
x"01700",-- 368
x"01b00",-- 432
x"01e00",-- 480
x"02300",-- 560
x"02700",-- 624
x"02b00",-- 688
x"02f00",-- 752
x"03100",-- 784
x"03500",-- 848
x"03900",-- 912
x"03c00",-- 960
x"03c00",-- 960
x"04000",-- 1024
x"04100",-- 1040
x"04100",-- 1040
x"04100",-- 1040
x"04100",-- 1040
x"03d00",-- 976
x"03900",-- 912
x"03800",-- 896
x"03700",-- 880
x"03300",-- 816
x"02e00",-- 736
x"02e00",-- 736
x"02c00",-- 704
x"02700",-- 624
x"02600",-- 608
x"02800",-- 640
x"02600",-- 608
x"02500",-- 592
x"02700",-- 624
x"02700",-- 624
x"02800",-- 640
x"02800",-- 640
x"02c00",-- 704
x"03000",-- 768
x"03400",-- 832
x"03700",-- 880
x"03a00",-- 928
x"04000",-- 1024
x"04600",-- 1120
x"04800",-- 1152
x"04900",-- 1168
x"04800",-- 1152
x"04300",-- 1072
x"03c00",-- 960
x"03700",-- 880
x"03300",-- 816
x"02800",-- 640
x"01d00",-- 464
x"01500",-- 336
x"00b00",-- 176
x"fff00",-- -16
x"ff600",-- -160
x"fec00",-- -320
x"fe400",-- -448
x"fdb00",-- -592
x"fd500",-- -688
x"fd600",-- -672
x"fd200",-- -736
x"fcf00",-- -784
x"fcc00",-- -832
x"fcc00",-- -832
x"fc800",-- -896
x"fc600",-- -928
x"fc600",-- -928
x"fc200",-- -992
x"fc200",-- -992
x"fbf00",-- -1040
x"fc100",-- -1008
x"fbf00",-- -1040
x"fba00",-- -1120
x"fb700",-- -1168
x"fb500",-- -1200
x"fb300",-- -1232
x"faf00",-- -1296
x"fb000",-- -1280
x"fb200",-- -1248
x"fae00",-- -1312
x"fb000",-- -1280
x"fb200",-- -1248
x"fb300",-- -1232
x"fb500",-- -1200
x"fb800",-- -1152
x"fbe00",-- -1056
x"fc200",-- -992
x"fc700",-- -912
x"fce00",-- -800
x"fd400",-- -704
x"fd700",-- -656
x"fdb00",-- -592
x"fe300",-- -464
x"fe900",-- -368
x"fed00",-- -304
x"ff200",-- -224
x"ff900",-- -112
x"ffd00",-- -48
x"00000",-- 0
x"00700",-- 112
x"00a00",-- 160
x"00d00",-- 208
x"01100",-- 272
x"01500",-- 336
x"01a00",-- 416
x"01b00",-- 432
x"01e00",-- 480
x"02000",-- 512
x"02100",-- 528
x"02200",-- 544
x"02400",-- 576
x"02700",-- 624
x"02600",-- 608
x"02600",-- 608
x"02800",-- 640
x"02700",-- 624
x"02600",-- 608
x"02500",-- 592
x"02500",-- 592
x"02200",-- 544
x"01f00",-- 496
x"01f00",-- 496
x"01e00",-- 480
x"01c00",-- 448
x"01800",-- 384
x"01700",-- 368
x"01500",-- 336
x"01100",-- 272
x"00f00",-- 240
x"00d00",-- 208
x"00c00",-- 192
x"00900",-- 144
x"00700",-- 112
x"00600",-- 96
x"00600",-- 96
x"00300",-- 48
x"00100",-- 16
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00700",-- 112
x"00a00",-- 160
x"00b00",-- 176
x"00d00",-- 208
x"01000",-- 256
x"01200",-- 288
x"01400",-- 320
x"01600",-- 352
x"01c00",-- 448
x"02100",-- 528
x"02300",-- 560
x"02500",-- 592
x"02a00",-- 672
x"02e00",-- 736
x"03200",-- 800
x"03700",-- 880
x"03800",-- 896
x"03900",-- 912
x"03500",-- 848
x"03100",-- 784
x"02f00",-- 752
x"02a00",-- 672
x"02600",-- 608
x"01f00",-- 496
x"01b00",-- 432
x"01300",-- 304
x"00b00",-- 176
x"00400",-- 64
x"ffc00",-- -64
x"ff500",-- -176
x"fef00",-- -272
x"fed00",-- -304
x"feb00",-- -336
x"fe800",-- -384
x"fe600",-- -416
x"fe600",-- -416
x"fe200",-- -480
x"fdf00",-- -528
x"fdf00",-- -528
x"fde00",-- -544
x"fdb00",-- -592
x"fda00",-- -608
x"fd900",-- -624
x"fd800",-- -640
x"fd800",-- -640
x"fd400",-- -704
x"fd000",-- -768
x"fce00",-- -800
x"fcb00",-- -848
x"fc800",-- -896
x"fc800",-- -896
x"fc700",-- -912
x"fc400",-- -960
x"fc200",-- -992
x"fc200",-- -992
x"fc100",-- -1008
x"fc200",-- -992
x"fc300",-- -976
x"fc600",-- -928
x"fc900",-- -880
x"fcc00",-- -832
x"fd100",-- -752
x"fd300",-- -720
x"fd800",-- -640
x"fda00",-- -608
x"fe100",-- -496
x"fe700",-- -400
x"fec00",-- -320
x"ff300",-- -208
x"ff700",-- -144
x"ffd00",-- -48
x"00100",-- 16
x"00800",-- 128
x"00d00",-- 208
x"01100",-- 272
x"01600",-- 352
x"01900",-- 400
x"01d00",-- 464
x"02100",-- 528
x"02400",-- 576
x"02600",-- 608
x"02800",-- 640
x"02900",-- 656
x"02a00",-- 672
x"02c00",-- 704
x"02c00",-- 704
x"02b00",-- 688
x"02b00",-- 688
x"02900",-- 656
x"02600",-- 608
x"02400",-- 576
x"02200",-- 544
x"01f00",-- 496
x"01b00",-- 432
x"01900",-- 400
x"01600",-- 352
x"01300",-- 304
x"01000",-- 256
x"00d00",-- 208
x"00a00",-- 160
x"00800",-- 128
x"00500",-- 80
x"00400",-- 64
x"00200",-- 32
x"00000",-- 0
x"ffe00",-- -32
x"ffc00",-- -64
x"ffa00",-- -96
x"ff800",-- -128
x"ff600",-- -160
x"ff400",-- -192
x"ff200",-- -224
x"ff100",-- -240
x"ff000",-- -256
x"fee00",-- -288
x"fed00",-- -304
x"fed00",-- -304
x"fec00",-- -320
x"fec00",-- -320
x"fee00",-- -288
x"fef00",-- -272
x"ff100",-- -240
x"ff200",-- -224
x"ff600",-- -160
x"ff800",-- -128
x"ffa00",-- -96
x"ffe00",-- -32
x"00300",-- 48
x"00600",-- 96
x"00900",-- 144
x"00e00",-- 224
x"01200",-- 288
x"01700",-- 368
x"01b00",-- 432
x"01f00",-- 496
x"02500",-- 592
x"02800",-- 640
x"02c00",-- 704
x"03000",-- 768
x"03300",-- 816
x"03400",-- 832
x"03400",-- 832
x"03300",-- 816
x"03100",-- 784
x"02f00",-- 752
x"02c00",-- 704
x"02800",-- 640
x"02400",-- 576
x"01e00",-- 480
x"01900",-- 400
x"01300",-- 304
x"00d00",-- 208
x"00800",-- 128
x"00400",-- 64
x"fff00",-- -16
x"ffb00",-- -80
x"ff800",-- -128
x"ff600",-- -160
x"ff400",-- -192
x"ff100",-- -240
x"fee00",-- -288
x"fec00",-- -320
x"fea00",-- -352
x"fe700",-- -400
x"fe600",-- -416
x"fe300",-- -464
x"fe000",-- -512
x"fde00",-- -544
x"fdb00",-- -592
x"fd800",-- -640
x"fd600",-- -672
x"fd300",-- -720
x"fd000",-- -768
x"fcf00",-- -784
x"fce00",-- -800
x"fcd00",-- -816
x"fcd00",-- -816
x"fcd00",-- -816
x"fcd00",-- -816
x"fce00",-- -800
x"fd100",-- -752
x"fd300",-- -720
x"fd600",-- -672
x"fda00",-- -608
x"fde00",-- -544
x"fe200",-- -480
x"fe600",-- -416
x"fea00",-- -352
x"fee00",-- -288
x"ff200",-- -224
x"ff600",-- -160
x"ffa00",-- -96
x"ffe00",-- -32
x"00100",-- 16
x"00400",-- 64
x"00600",-- 96
x"00900",-- 144
x"00b00",-- 176
x"00d00",-- 208
x"00f00",-- 240
x"01100",-- 272
x"01300",-- 304
x"01400",-- 320
x"01500",-- 336
x"01500",-- 336
x"01600",-- 352
x"01500",-- 336
x"01500",-- 336
x"01600",-- 352
x"01500",-- 336
x"01600",-- 352
x"01500",-- 336
x"01500",-- 336
x"01400",-- 320
x"01300",-- 304
x"01300",-- 304
x"01200",-- 288
x"01200",-- 288
x"01000",-- 256
x"01000",-- 256
x"01000",-- 256
x"00e00",-- 224
x"00c00",-- 192
x"00b00",-- 176
x"00900",-- 144
x"00900",-- 144
x"00600",-- 96
x"00500",-- 80
x"00300",-- 48
x"00200",-- 32
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00300",-- 48
x"00500",-- 80
x"00600",-- 96
x"00800",-- 128
x"00a00",-- 160
x"00c00",-- 192
x"00f00",-- 240
x"01200",-- 288
x"01500",-- 336
x"01700",-- 368
x"01b00",-- 432
x"01e00",-- 480
x"02000",-- 512
x"02300",-- 560
x"02300",-- 560
x"02400",-- 576
x"02300",-- 560
x"02200",-- 544
x"02100",-- 528
x"01f00",-- 496
x"01c00",-- 448
x"01800",-- 384
x"01600",-- 352
x"01000",-- 256
x"00c00",-- 192
x"00800",-- 128
x"00400",-- 64
x"00000",-- 0
x"ffc00",-- -64
x"ffa00",-- -96
x"ff700",-- -144
x"ff500",-- -176
x"ff200",-- -224
x"ff100",-- -240
x"fef00",-- -272
x"fec00",-- -320
x"feb00",-- -336
x"fea00",-- -352
x"fe800",-- -384
x"fe600",-- -416
x"fe500",-- -432
x"fe400",-- -448
x"fe300",-- -464
x"fe000",-- -512
x"fdf00",-- -528
x"fdf00",-- -528
x"fdc00",-- -576
x"fdc00",-- -576
x"fdb00",-- -592
x"fdb00",-- -592
x"fd900",-- -624
x"fda00",-- -608
x"fdb00",-- -592
x"fdb00",-- -592
x"fdc00",-- -576
x"fdd00",-- -560
x"fdf00",-- -528
x"fe100",-- -496
x"fe300",-- -464
x"fe600",-- -416
x"fe800",-- -384
x"fea00",-- -352
x"fec00",-- -320
x"ff000",-- -256
x"ff200",-- -224
x"ff400",-- -192
x"ff700",-- -144
x"ff800",-- -128
x"ffa00",-- -96
x"ffc00",-- -64
x"ffe00",-- -32
x"00000",-- 0
x"00200",-- 32
x"00300",-- 48
x"00600",-- 96
x"00900",-- 144
x"00900",-- 144
x"00c00",-- 192
x"00e00",-- 224
x"00f00",-- 240
x"01000",-- 256
x"01200",-- 288
x"01300",-- 304
x"01300",-- 304
x"01400",-- 320
x"01400",-- 320
x"01300",-- 304
x"01300",-- 304
x"01200",-- 288
x"01200",-- 288
x"01200",-- 288
x"01200",-- 288
x"01100",-- 272
x"01100",-- 272
x"01000",-- 256
x"00f00",-- 240
x"00f00",-- 240
x"00e00",-- 224
x"00d00",-- 208
x"00d00",-- 208
x"00d00",-- 208
x"00b00",-- 176
x"00b00",-- 176
x"00900",-- 144
x"00900",-- 144
x"00800",-- 128
x"00700",-- 112
x"00700",-- 112
x"00500",-- 80
x"00500",-- 80
x"00500",-- 80
x"00500",-- 80
x"00400",-- 64
x"00300",-- 48
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00500",-- 80
x"00600",-- 96
x"00600",-- 96
x"00800",-- 128
x"00900",-- 144
x"00b00",-- 176
x"00c00",-- 192
x"00e00",-- 224
x"01000",-- 256
x"01100",-- 272
x"01300",-- 304
x"01500",-- 336
x"01800",-- 384
x"01800",-- 384
x"01900",-- 400
x"01b00",-- 432
x"01c00",-- 448
x"01b00",-- 432
x"01b00",-- 432
x"01a00",-- 416
x"01800",-- 384
x"01600",-- 352
x"01400",-- 320
x"01100",-- 272
x"00f00",-- 240
x"00b00",-- 176
x"00800",-- 128
x"00500",-- 80
x"00000",-- 0
x"ffd00",-- -48
x"ffb00",-- -80
x"ff700",-- -144
x"ff300",-- -208
x"ff200",-- -224
x"ff000",-- -256
x"fed00",-- -304
x"fec00",-- -320
x"fea00",-- -352
x"fe800",-- -384
x"fe500",-- -432
x"fe400",-- -448
x"fe300",-- -464
x"fe200",-- -480
x"fe000",-- -512
x"fdf00",-- -528
x"fdf00",-- -528
x"fdd00",-- -560
x"fdc00",-- -576
x"fdc00",-- -576
x"fdb00",-- -592
x"fda00",-- -608
x"fdb00",-- -592
x"fdb00",-- -592
x"fdc00",-- -576
x"fdd00",-- -560
x"fdd00",-- -560
x"fe000",-- -512
x"fe200",-- -480
x"fe300",-- -464
x"fe600",-- -416
x"fe900",-- -368
x"fec00",-- -320
x"fee00",-- -288
x"ff100",-- -240
x"ff400",-- -192
x"ff700",-- -144
x"ff900",-- -112
x"ffd00",-- -48
x"00000",-- 0
x"00300",-- 48
x"00500",-- 80
x"00800",-- 128
x"00a00",-- 160
x"00c00",-- 192
x"00f00",-- 240
x"01100",-- 272
x"01300",-- 304
x"01400",-- 320
x"01500",-- 336
x"01700",-- 368
x"01800",-- 384
x"01800",-- 384
x"01900",-- 400
x"01b00",-- 432
x"01a00",-- 416
x"01b00",-- 432
x"01b00",-- 432
x"01a00",-- 416
x"01900",-- 400
x"01900",-- 400
x"01800",-- 384
x"01700",-- 368
x"01600",-- 352
x"01500",-- 336
x"01400",-- 320
x"01200",-- 288
x"01100",-- 272
x"00f00",-- 240
x"00e00",-- 224
x"00c00",-- 192
x"00a00",-- 160
x"00900",-- 144
x"00800",-- 128
x"00600",-- 96
x"00500",-- 80
x"00300",-- 48
x"00200",-- 32
x"00000",-- 0
x"fff00",-- -16
x"ffd00",-- -48
x"ffc00",-- -64
x"ffc00",-- -64
x"ffb00",-- -80
x"ffb00",-- -80
x"ff900",-- -112
x"ff900",-- -112
x"ff900",-- -112
x"ff800",-- -128
x"ff900",-- -112
x"ff900",-- -112
x"ff900",-- -112
x"ff900",-- -112
x"ffa00",-- -96
x"ffb00",-- -80
x"ffb00",-- -80
x"ffb00",-- -80
x"ffc00",-- -64
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00300",-- 48
x"00300",-- 48
x"00300",-- 48
x"00200",-- 32
x"00300",-- 48
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffd00",-- -48
x"ffc00",-- -64
x"ffc00",-- -64
x"ffb00",-- -80
x"ff900",-- -112
x"ffa00",-- -96
x"ff900",-- -112
x"ff800",-- -128
x"ff700",-- -144
x"ff700",-- -144
x"ff700",-- -144
x"ff600",-- -160
x"ff600",-- -160
x"ff600",-- -160
x"ff500",-- -176
x"ff400",-- -192
x"ff400",-- -192
x"ff500",-- -176
x"ff400",-- -192
x"ff400",-- -192
x"ff400",-- -192
x"ff500",-- -176
x"ff500",-- -176
x"ff500",-- -176
x"ff700",-- -144
x"ff700",-- -144
x"ff700",-- -144
x"ff700",-- -144
x"ff900",-- -112
x"ffa00",-- -96
x"ffa00",-- -96
x"ffb00",-- -80
x"ffc00",-- -64
x"ffd00",-- -48
x"ffd00",-- -48
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"00300",-- 48
x"00500",-- 80
x"00500",-- 80
x"00600",-- 96
x"00600",-- 96
x"00800",-- 128
x"00800",-- 128
x"00900",-- 144
x"00a00",-- 160
x"00a00",-- 160
x"00a00",-- 160
x"00a00",-- 160
x"00b00",-- 176
x"00b00",-- 176
x"00b00",-- 176
x"00a00",-- 160
x"00b00",-- 176
x"00a00",-- 160
x"00900",-- 144
x"00a00",-- 160
x"00900",-- 144
x"00900",-- 144
x"00800",-- 128
x"00800",-- 128
x"00700",-- 112
x"00700",-- 112
x"00600",-- 96
x"00500",-- 80
x"00400",-- 64
x"00400",-- 64
x"00300",-- 48
x"00300",-- 48
x"00200",-- 32
x"00100",-- 16
x"00000",-- 0
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffc00",-- -64
x"ffc00",-- -64
x"ffb00",-- -80
x"ffb00",-- -80
x"ffa00",-- -96
x"ffa00",-- -96
x"ffa00",-- -96
x"ff900",-- -112
x"ff900",-- -112
x"ff800",-- -128
x"ff800",-- -128
x"ff900",-- -112
x"ff800",-- -128
x"ff800",-- -128
x"ff800",-- -128
x"ff800",-- -128
x"ff800",-- -128
x"ff900",-- -112
x"ff900",-- -112
x"ffa00",-- -96
x"ffa00",-- -96
x"ffb00",-- -80
x"ffb00",-- -80
x"ffc00",-- -64
x"ffc00",-- -64
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00300",-- 48
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00500",-- 80
x"00300",-- 48
x"00400",-- 64
x"00500",-- 80
x"00400",-- 64
x"00400",-- 64
x"00500",-- 80
x"00400",-- 64
x"00400",-- 64
x"00500",-- 80
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00300",-- 48
x"00300",-- 48
x"00300",-- 48
x"00300",-- 48
x"00300",-- 48
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffd00",-- -48
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffc00",-- -64
x"ffc00",-- -64
x"ffd00",-- -48
x"ffc00",-- -64
x"ffc00",-- -64
x"ffd00",-- -48
x"ffc00",-- -64
x"ffc00",-- -64
x"ffc00",-- -64
x"ffc00",-- -64
x"ffc00",-- -64
x"ffc00",-- -64
x"ffc00",-- -64
x"ffd00",-- -48
x"ffd00",-- -48
x"ffc00",-- -64
x"ffd00",-- -48
x"ffd00",-- -48
x"ffd00",-- -48
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00300",-- 48
x"00300",-- 48
x"00300",-- 48
x"00300",-- 48
x"00300",-- 48
x"00300",-- 48
x"00300",-- 48
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00500",-- 80
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00500",-- 80
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00300",-- 48
x"00400",-- 64
x"00400",-- 64
x"00400",-- 64
x"00300",-- 48
x"00300",-- 48
x"00300",-- 48
x"00300",-- 48
x"00200",-- 32
x"00300",-- 48
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00100",-- 16
x"00200",-- 32
x"00200",-- 32
x"00100",-- 16
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00100",-- 16
x"00100",-- 16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff00",-- -16
x"fff00",-- -16
x"fff00",-- -16
x"ffe00",-- -32
x"ffe00",-- -32
x"ffc00",-- -64
x"ffc00",-- -64
x"ff800",-- -128
x"ff500",-- -176
x"fed00",-- -304
x"fe600",-- -416
x"fc200",-- -992
x"f7900",-- -2160
x"fe700",-- -400
x"05c00",-- 1472
x"01e00",-- 480
x"00400",-- 64
x"00800",-- 128
x"01100",-- 272
x"00f00",-- 240
x"00c00",-- 192
x"00c00",-- 192
x"ff700",-- -144
x"00600",-- 96
x"01100",-- 272
x"01100",-- 272
x"01b00",-- 432
x"02600",-- 608
x"02800",-- 640
x"01b00",-- 432
x"00600",-- 96
x"00800",-- 128
x"00a00",-- 160
x"fef00",-- -272
x"00800",-- 128
x"fff00",-- -16
x"fde00",-- -544
x"ff900",-- -112
x"ff900",-- -112
x"ff600",-- -160
x"ff800",-- -128
x"ff000",-- -256
x"ff100",-- -240
x"00500",-- 80
x"00100",-- 16
x"00000",-- 0
x"01000",-- 256
x"00300",-- 48
x"fdf00",-- -528
x"ffb00",-- -80
x"01100",-- 272
x"fe900",-- -368
x"ff700",-- -144
x"ffe00",-- -32
x"00500",-- 80
x"00300",-- 48
x"ff200",-- -224
x"01000",-- 256
x"00900",-- 144
x"ff000",-- -256
x"00700",-- 112
x"01000",-- 256
x"00400",-- 64
x"00900",-- 144
x"00a00",-- 160
x"ffd00",-- -48
x"ffc00",-- -64
x"01100",-- 272
x"ffe00",-- -32
x"ff200",-- -224
x"01800",-- 384
x"ff500",-- -176
x"00900",-- 144
x"00000",-- 0
x"fe700",-- -400
x"00e00",-- 224
x"ff200",-- -224
x"fda00",-- -608
x"00400",-- 64
x"00700",-- 112
x"fbc00",-- -1088
x"fe100",-- -496
x"ff700",-- -144
x"fd000",-- -768
x"01900",-- 400
x"ffb00",-- -80
x"fee00",-- -288
x"02a00",-- 672
x"ff400",-- -192
x"01d00",-- 464
x"01200",-- 288
x"ff100",-- -240
x"01600",-- 352
x"02f00",-- 752
x"00a00",-- 160
x"01c00",-- 448
x"fd700",-- -656
x"fa700",-- -1424
x"03900",-- 912
x"fe700",-- -400
x"ffa00",-- -96
x"06200",-- 1568
x"f9f00",-- -1552
x"01a00",-- 416
x"07000",-- 1792
x"f9500",-- -1712
x"05400",-- 1344
x"03100",-- 784
x"fa400",-- -1472
x"04500",-- 1104
x"01400",-- 320
x"fec00",-- -320
x"00c00",-- 192
x"04b00",-- 1200
x"00e00",-- 224
x"01a00",-- 416
x"07200",-- 1824
x"fa800",-- -1408
x"03100",-- 784
x"02700",-- 624
x"fc000",-- -1024
x"04700",-- 1136
x"fab00",-- -1360
x"01d00",-- 464
x"00700",-- 112
x"fbc00",-- -1088
x"02100",-- 528
x"fc400",-- -960
x"f7100",-- -2288
x"fe400",-- -448
x"0a300",-- 2608
x"fd100",-- -752
x"00600",-- 96
x"03c00",-- 960
x"f8d00",-- -1840
x"fed00",-- -304
x"04200",-- 1056
x"faa00",-- -1376
x"fd200",-- -736
x"04d00",-- 1232
x"fd900",-- -624
x"02500",-- 592
x"02300",-- 560
x"feb00",-- -336
x"06700",-- 1648
x"02200",-- 544
x"fc500",-- -944
x"04b00",-- 1200
x"fcd00",-- -816
x"fea00",-- -352
x"03c00",-- 960
x"00a00",-- 160
x"00800",-- 128
x"ffa00",-- -96
x"04900",-- 1168
x"fc000",-- -1024
x"01a00",-- 416
x"fe400",-- -448
x"f8700",-- -1936
x"00400",-- 64
x"fab00",-- -1360
x"00200",-- 32
x"ff000",-- -256
x"fa100",-- -1520
x"00b00",-- 176
x"fe900",-- -368
x"ffa00",-- -96
x"05a00",-- 1440
x"fee00",-- -288
x"03e00",-- 992
x"04c00",-- 1216
x"fbf00",-- -1040
x"00f00",-- 240
x"03200",-- 800
x"faf00",-- -1296
x"ffd00",-- -48
x"02b00",-- 688
x"fab00",-- -1360
x"04f00",-- 1264
x"fce00",-- -800
x"03800",-- 896
x"07f00",-- 2032
x"f9b00",-- -1616
x"03f00",-- 1008
x"fed00",-- -304
x"fdb00",-- -592
x"00100",-- 16
x"ffc00",-- -64
x"fe200",-- -480
x"ff900",-- -112
x"01400",-- 320
x"fd000",-- -768
x"07000",-- 1792
x"fcc00",-- -832
x"00e00",-- 224
x"03000",-- 768
x"fcf00",-- -784
x"03400",-- 832
x"ffb00",-- -80
x"fee00",-- -288
x"01500",-- 336
x"fd700",-- -656
x"fd300",-- -720
x"03000",-- 768
x"ff200",-- -224
x"fa200",-- -1504
x"06500",-- 1616
x"00a00",-- 160
x"fb400",-- -1216
x"07500",-- 1872
x"00200",-- 32
x"fd100",-- -752
x"04300",-- 1072
x"ff500",-- -176
x"00a00",-- 160
x"02a00",-- 672
x"fcc00",-- -832
x"02300",-- 560
x"02d00",-- 720
x"fb000",-- -1280
x"01500",-- 336
x"04500",-- 1104
x"fa000",-- -1536
x"02400",-- 576
x"03c00",-- 960
x"fa700",-- -1424
x"04f00",-- 1264
x"ff600",-- -160
x"fb600",-- -1184
x"07100",-- 1808
x"fc400",-- -960
x"fe800",-- -384
x"05900",-- 1424
x"fb600",-- -1184
x"01000",-- 256
x"00b00",-- 176
x"ff100",-- -240
x"00f00",-- 240
x"fe000",-- -512
x"03100",-- 784
x"fe600",-- -416
x"01a00",-- 416
x"fec00",-- -320
x"ffb00",-- -80
x"01f00",-- 496
x"fc100",-- -1008
x"06300",-- 1584
x"f9900",-- -1648
x"00d00",-- 208
x"05800",-- 1408
x"f6b00",-- -2384
x"03c00",-- 960
x"03300",-- 816
x"f9f00",-- -1552
x"00200",-- 32
x"06100",-- 1552
x"fc300",-- -976
x"ff200",-- -224
x"02f00",-- 752
x"ff000",-- -256
x"fe200",-- -480
x"ffa00",-- -96
x"02a00",-- 672
x"fd600",-- -672
x"ffc00",-- -64
x"03300",-- 816
x"fcd00",-- -816
x"ff000",-- -256
x"02100",-- 528
x"fea00",-- -352
x"fe300",-- -464
x"02000",-- 512
x"00800",-- 128
x"fb700",-- -1168
x"01e00",-- 480
x"00400",-- 64
x"fcf00",-- -784
x"03f00",-- 1008
x"ffd00",-- -48
x"fcf00",-- -784
x"01500",-- 336
x"00600",-- 96
x"00e00",-- 224
x"fca00",-- -864
x"ffb00",-- -80
x"02000",-- 512
x"01000",-- 256
x"fd900",-- -624
x"00d00",-- 208
x"01100",-- 272
x"f9900",-- -1648
x"05700",-- 1392
x"01800",-- 384
x"fbb00",-- -1104
x"02900",-- 656
x"00600",-- 96
x"fe200",-- -480
x"00b00",-- 176
x"01b00",-- 432
x"fd800",-- -640
x"00700",-- 112
x"ff200",-- -224
x"ffa00",-- -96
x"01900",-- 400
x"fed00",-- -304
x"01500",-- 336
x"00200",-- 32
x"fc700",-- -912
x"02f00",-- 752
x"ff700",-- -144
x"fec00",-- -320
x"03c00",-- 960
x"fae00",-- -1312
x"00b00",-- 176
x"02a00",-- 672
x"fd100",-- -752
x"fd200",-- -736
x"04100",-- 1040
x"fda00",-- -608
x"fd000",-- -768
x"09d00",-- 2512
x"f9a00",-- -1632
x"fe600",-- -416
x"03f00",-- 1008
x"fef00",-- -272
x"02600",-- 608
x"fbf00",-- -1040
x"02800",-- 640
x"fe400",-- -448
x"fdc00",-- -576
x"fff00",-- -16
x"fd400",-- -704
x"03200",-- 800
x"00400",-- 64
x"fe300",-- -464
x"02b00",-- 688
x"ff700",-- -144
x"ff200",-- -224
x"01500",-- 336
x"01400",-- 320
x"01900",-- 400
x"fdb00",-- -592
x"01600",-- 352
x"00e00",-- 224
x"fc500",-- -944
x"00800",-- 128
x"01200",-- 288
x"01c00",-- 448
x"fd800",-- -640
x"fda00",-- -608
x"03d00",-- 976
x"fdc00",-- -576
x"fa500",-- -1456
x"03400",-- 832
x"fda00",-- -608
x"fd000",-- -768
x"00b00",-- 176
x"ff400",-- -192
x"00200",-- 32
x"fda00",-- -608
x"04200",-- 1056
x"00500",-- 80
x"fe900",-- -368
x"02f00",-- 752
x"00500",-- 80
x"02a00",-- 672
x"01b00",-- 432
x"fdb00",-- -592
x"02a00",-- 672
x"06b00",-- 1712
x"fd300",-- -720
x"ff900",-- -112
x"04700",-- 1136
x"00300",-- 48
x"fc200",-- -992
x"04900",-- 1168
x"00d00",-- 208
x"f9200",-- -1760
x"06600",-- 1632
x"fa800",-- -1408
x"05400",-- 1344
x"fe100",-- -496
x"f6100",-- -2544
x"0cc00",-- 3264
x"f5100",-- -2800
x"01700",-- 368
x"04000",-- 1024
x"f9000",-- -1792
x"05300",-- 1328
x"fcd00",-- -816
x"03300",-- 816
x"00000",-- 0
x"00700",-- 112
x"03900",-- 912
x"f8400",-- -1984
x"0b500",-- 2896
x"00400",-- 64
x"fca00",-- -864
x"02900",-- 656
x"fd900",-- -624
x"08e00",-- 2272
x"f7900",-- -2160
x"07300",-- 1840
x"fcb00",-- -848
x"fe800",-- -384
x"0b500",-- 2896
x"f1700",-- -3728
x"0b400",-- 2880
x"00500",-- 80
x"f3a00",-- -3168
x"0db00",-- 3504
x"fd400",-- -704
x"fa500",-- -1456
x"04a00",-- 1184
x"fc200",-- -992
x"00c00",-- 192
x"fff00",-- -16
x"01000",-- 256
x"fe900",-- -368
x"fd600",-- -672
x"fef00",-- -272
x"02a00",-- 672
x"04f00",-- 1264
x"f5d00",-- -2608
x"02700",-- 624
x"07400",-- 1856
x"f8900",-- -1904
x"04a00",-- 1184
x"03800",-- 896
x"f9600",-- -1696
x"00800",-- 128
x"05c00",-- 1472
x"ff600",-- -160
x"f9600",-- -1696
x"08400",-- 2112
x"ff000",-- -256
x"f9c00",-- -1600
x"0b000",-- 2816
x"f8700",-- -1936
x"00e00",-- 224
x"03400",-- 832
x"f7200",-- -2272
x"0a500",-- 2640
x"fef00",-- -272
x"f7e00",-- -2080
x"03800",-- 896
x"ff900",-- -112
x"fe700",-- -400
x"00600",-- 96
x"ff800",-- -128
x"00000",-- 0
x"02000",-- 512
x"fc300",-- -976
x"01500",-- 336
x"02200",-- 544
x"fc400",-- -960
x"feb00",-- -336
x"03f00",-- 1008
x"fe800",-- -384
x"fe500",-- -432
x"01600",-- 352
x"fdb00",-- -592
x"02500",-- 592
x"fcb00",-- -848
x"02400",-- 576
x"00700",-- 112
x"fb900",-- -1136
x"07d00",-- 2000
x"fab00",-- -1360
x"ff900",-- -112
x"04f00",-- 1264
x"f7a00",-- -2144
x"04500",-- 1104
x"03500",-- 848
x"fa100",-- -1520
x"02600",-- 608
x"00600",-- 96
x"fdf00",-- -528
x"00c00",-- 192
x"01200",-- 288
x"ff200",-- -224
x"ff700",-- -144
x"00700",-- 112
x"fd600",-- -672
x"03700",-- 880
x"00400",-- 64
x"fc700",-- -912
x"02500",-- 592
x"02100",-- 528
x"fff00",-- -16
x"00b00",-- 176
x"00c00",-- 192
x"fd000",-- -768
x"03e00",-- 992
x"00900",-- 144
x"f9b00",-- -1616
x"05a00",-- 1440
x"ffa00",-- -96
x"fbb00",-- -1104
x"04f00",-- 1264
x"fe500",-- -432
x"ffc00",-- -64
x"01d00",-- 464
x"fe400",-- -448
x"ffe00",-- -32
x"02a00",-- 672
x"00900",-- 144
x"fd800",-- -640
x"01600",-- 352
x"ffe00",-- -32
x"ffa00",-- -96
x"00000",-- 0
x"fe300",-- -464
x"feb00",-- -336
x"02300",-- 560
x"02c00",-- 704
x"fe400",-- -448
x"fcb00",-- -848
x"03500",-- 848
x"01800",-- 384
x"fd400",-- -704
x"03600",-- 864
x"fed00",-- -304
x"fe000",-- -512
x"01100",-- 272
x"00d00",-- 208
x"01700",-- 368
x"fe300",-- -464
x"00300",-- 48
x"fe700",-- -400
x"00e00",-- 224
x"02600",-- 608
x"fbe00",-- -1056
x"02f00",-- 752
x"fdd00",-- -560
x"00b00",-- 176
x"04200",-- 1056
x"fc900",-- -880
x"ff700",-- -144
x"01700",-- 368
x"fe400",-- -448
x"04400",-- 1088
x"fdd00",-- -560
x"00900",-- 144
x"01b00",-- 432
x"f9b00",-- -1616
x"07300",-- 1840
x"00e00",-- 224
x"fad00",-- -1328
x"02600",-- 608
x"01400",-- 320
x"ff300",-- -208
x"00600",-- 96
x"01100",-- 272
x"fd200",-- -736
x"03000",-- 768
x"feb00",-- -336
x"00200",-- 32
x"04600",-- 1120
x"fc500",-- -944
x"fe600",-- -416
x"03100",-- 784
x"00500",-- 80
x"fff00",-- -16
x"ff200",-- -224
x"fc700",-- -912
x"02500",-- 592
x"01300",-- 304
x"ff400",-- -192
x"00d00",-- 208
x"fe100",-- -496
x"00200",-- 32
x"03f00",-- 1008
x"fda00",-- -608
x"fe600",-- -416
x"02a00",-- 672
x"fdc00",-- -576
x"fe500",-- -432
x"02d00",-- 720
x"ff500",-- -176
x"00200",-- 32
x"00c00",-- 192
x"fc600",-- -928
x"02200",-- 544
x"03f00",-- 1008
x"fc900",-- -880
x"ff200",-- -224
x"02500",-- 592
x"00a00",-- 160
x"02900",-- 656
x"ff100",-- -240
x"fcf00",-- -784
x"03200",-- 800
x"01200",-- 288
x"ff900",-- -112
x"01d00",-- 464
x"fed00",-- -304
x"fd700",-- -656
x"00400",-- 64
x"01700",-- 368
x"01000",-- 256
x"fe000",-- -512
x"fd900",-- -624
x"02500",-- 592
x"00c00",-- 192
x"fea00",-- -352
x"ff500",-- -176
x"ff300",-- -208
x"01700",-- 368
x"ff100",-- -240
x"fde00",-- -544
x"02600",-- 608
x"00700",-- 112
x"fe500",-- -432
x"01e00",-- 480
x"02a00",-- 672
x"fe900",-- -368
x"ff200",-- -224
x"01200",-- 288
x"02500",-- 592
x"fff00",-- -16
x"ffa00",-- -96
x"00500",-- 80
x"fe400",-- -448
x"00200",-- 32
x"ffa00",-- -96
x"fee00",-- -288
x"02a00",-- 672
x"01100",-- 272
x"fe300",-- -464
x"00500",-- 80
x"00700",-- 112
x"fe800",-- -384
x"00f00",-- 240
x"01100",-- 272
x"fe500",-- -432
x"00a00",-- 160
x"fd800",-- -640
x"ff900",-- -112
x"03e00",-- 992
x"fb500",-- -1200
x"ffa00",-- -96
x"03100",-- 784
x"fe500",-- -432
x"ff300",-- -208
x"02300",-- 560
x"00300",-- 48
x"feb00",-- -336
x"00c00",-- 192
x"fe500",-- -432
x"02b00",-- 688
x"00c00",-- 192
x"fca00",-- -864
x"03900",-- 912
x"00d00",-- 208
x"fc700",-- -912
x"00900",-- 144
x"01200",-- 288
x"fec00",-- -320
x"00200",-- 32
x"00100",-- 16
x"ff200",-- -224
x"ffe00",-- -32
x"fe100",-- -496
x"ffa00",-- -96
x"02500",-- 592
x"ff100",-- -240
x"ff000",-- -256
x"01600",-- 352
x"ff500",-- -176
x"fe300",-- -464
x"01d00",-- 464
x"01900",-- 400
x"ff200",-- -224
x"ff000",-- -256
x"ff200",-- -224
x"02300",-- 560
x"ffe00",-- -32
x"fe800",-- -384
x"00a00",-- 160
x"01300",-- 304
x"fdd00",-- -560
x"00400",-- 64
x"01b00",-- 432
x"ff300",-- -208
x"fed00",-- -304
x"00300",-- 48
x"02100",-- 528
x"ffe00",-- -32
x"fed00",-- -304
x"00100",-- 16
x"01500",-- 336
x"00200",-- 32
x"00b00",-- 176
x"00d00",-- 208
x"ffb00",-- -80
x"ff100",-- -240
x"ffc00",-- -64
x"00e00",-- 224
x"01100",-- 272
x"ff000",-- -256
x"ff500",-- -176
x"01f00",-- 496
x"00400",-- 64
x"fed00",-- -304
x"01200",-- 288
x"ff300",-- -208
x"fe600",-- -416
x"01600",-- 352
x"fe300",-- -464
x"fe600",-- -416
x"00800",-- 128
x"ffa00",-- -96
x"01400",-- 320
x"fff00",-- -16
x"ffb00",-- -80
x"fe500",-- -432
x"ffc00",-- -64
x"01700",-- 368
x"00400",-- 64
x"00000",-- 0
x"00200",-- 32
x"ff800",-- -128
x"ffd00",-- -48
x"01e00",-- 480
x"00800",-- 128
x"fee00",-- -288
x"00d00",-- 208
x"00900",-- 144
x"00900",-- 144
x"01400",-- 320
x"ff900",-- -112
x"00000",-- 0
x"00000",-- 0
x"ffc00",-- -64
x"00000",-- 0
x"fe000",-- -512
x"fe300",-- -464
x"fe500",-- -432
x"00600",-- 96
x"01600",-- 352
x"fdb00",-- -592
x"fea00",-- -352
x"00600",-- 96
x"ffe00",-- -32
x"00600",-- 96
x"00100",-- 16
x"ff500",-- -176
x"ff800",-- -128
x"01e00",-- 480
x"00c00",-- 192
x"fe900",-- -368
x"ffc00",-- -64
x"01700",-- 368
x"00f00",-- 240
x"ffb00",-- -80
x"00b00",-- 176
x"00400",-- 64
x"ff400",-- -192
x"ff400",-- -192
x"00b00",-- 176
x"ffa00",-- -96
x"fef00",-- -272
x"01100",-- 272
x"01500",-- 336
x"ffd00",-- -48
x"fe800",-- -384
x"fe600",-- -416
x"00600",-- 96
x"00600",-- 96
x"ff000",-- -256
x"01d00",-- 464
x"ffb00",-- -80
x"fe000",-- -512
x"00c00",-- 192
x"00d00",-- 208
x"00a00",-- 160
x"01f00",-- 496
x"00300",-- 48
x"ff500",-- -176
x"00a00",-- 160
x"00f00",-- 240
x"01400",-- 320
x"ff800",-- -128
x"ff800",-- -128
x"00600",-- 96
x"00900",-- 144
x"ffc00",-- -64
x"00500",-- 80
x"ffd00",-- -48
x"fe100",-- -496
x"00200",-- 32
x"00e00",-- 224
x"ff700",-- -144
x"00100",-- 16
x"fff00",-- -16
x"ff600",-- -160
x"00600",-- 96
x"00a00",-- 160
x"ffe00",-- -32
x"ff800",-- -128
x"ff800",-- -128
x"ff200",-- -224
x"01000",-- 256
x"00f00",-- 240
x"ff300",-- -208
x"00900",-- 144
x"01000",-- 256
x"ff800",-- -128
x"ffb00",-- -80
x"00b00",-- 176
x"00300",-- 48
x"ff900",-- -112
x"ffa00",-- -96
x"01100",-- 272
x"00300",-- 48
x"fec00",-- -320
x"00800",-- 128
x"ff500",-- -176
x"ffe00",-- -32
x"01900",-- 400
x"00900",-- 144
x"00100",-- 16
x"00d00",-- 208
x"01200",-- 288
x"ff000",-- -256
x"ff500",-- -176
x"01300",-- 304
x"00900",-- 144
x"ff700",-- -144
x"fe700",-- -400
x"ff100",-- -240
x"00000",-- 0
x"00e00",-- 224
x"00800",-- 128
x"fdf00",-- -528
x"fe100",-- -496
x"00900",-- 144
x"01300",-- 304
x"00200",-- 32
x"ff800",-- -128
x"ff100",-- -240
x"00300",-- 48
x"02a00",-- 672
x"02400",-- 576
x"fef00",-- -272
x"fe200",-- -480
x"ff500",-- -176
x"01d00",-- 464
x"02a00",-- 672
x"00000",-- 0
x"fe700",-- -400
x"fed00",-- -304
x"00100",-- 16
x"00a00",-- 160
x"ffd00",-- -48
x"fe200",-- -480
x"fdd00",-- -560
x"ff000",-- -256
x"00900",-- 144
x"00b00",-- 176
x"fec00",-- -320
x"fd400",-- -704
x"fe100",-- -496
x"ff100",-- -240
x"00a00",-- 160
x"01b00",-- 432
x"ffa00",-- -96
x"ff200",-- -224
x"ff800",-- -128
x"00000",-- 0
x"ff600",-- -160
x"00100",-- 16
x"01400",-- 320
x"ffa00",-- -96
x"ff800",-- -128
x"00400",-- 64
x"00500",-- 80
x"ffc00",-- -64
x"ff900",-- -112
x"01700",-- 368
x"00800",-- 128
x"fc900",-- -880
x"fe500",-- -432
x"00a00",-- 160
x"00700",-- 112
x"00400",-- 64
x"ff000",-- -256
x"ffe00",-- -32
x"00300",-- 48
x"00e00",-- 224
x"01600",-- 352
x"00c00",-- 192
x"00700",-- 112
x"ff200",-- -224
x"fff00",-- -16
x"01e00",-- 480
x"01a00",-- 416
x"ffa00",-- -96
x"00400",-- 64
x"01700",-- 368
x"00200",-- 32
x"ff500",-- -176
x"00900",-- 144
x"00200",-- 32
x"ff100",-- -240
x"ffe00",-- -32
x"00600",-- 96
x"01400",-- 320
x"00100",-- 16
x"fec00",-- -320
x"ff100",-- -240
x"fed00",-- -304
x"ffd00",-- -48
x"01b00",-- 432
x"01400",-- 320
x"ff800",-- -128
x"00000",-- 0
x"01c00",-- 448
x"01600",-- 352
x"ffd00",-- -48
x"00000",-- 0
x"00300",-- 48
x"01100",-- 272
x"01400",-- 320
x"00400",-- 64
x"ff800",-- -128
x"ff500",-- -176
x"ff300",-- -208
x"ffd00",-- -48
x"00a00",-- 160
x"ff600",-- -160
x"fe700",-- -400
x"ff900",-- -112
x"00300",-- 48
x"ffe00",-- -32
x"ff000",-- -256
x"fea00",-- -352
x"ff500",-- -176
x"ffd00",-- -48
x"01700",-- 368
x"02100",-- 528
x"00d00",-- 208
x"ffe00",-- -32
x"ff400",-- -192
x"00000",-- 0
x"00100",-- 16
x"00200",-- 32
x"01300",-- 304
x"01000",-- 256
x"ffc00",-- -64
x"ffb00",-- -80
x"00900",-- 144
x"00900",-- 144
x"00800",-- 128
x"00400",-- 64
x"ff700",-- -144
x"ffd00",-- -48
x"00800",-- 128
x"00b00",-- 176
x"00400",-- 64
x"ffe00",-- -32
x"00100",-- 16
x"00900",-- 144
x"00300",-- 48
x"ff500",-- -176
x"ff400",-- -192
x"ff300",-- -208
x"ffd00",-- -48
x"00f00",-- 240
x"01900",-- 400
x"ff700",-- -144
x"fdd00",-- -560
x"ff700",-- -144
x"00400",-- 64
x"01000",-- 256
x"00a00",-- 160
x"fec00",-- -320
x"fe800",-- -384
x"ffe00",-- -32
x"ffc00",-- -64
x"ff800",-- -128
x"00000",-- 0
x"fef00",-- -272
x"ff200",-- -224
x"01600",-- 352
x"00e00",-- 224
x"fe900",-- -368
x"fe900",-- -368
x"ffd00",-- -48
x"00200",-- 32
x"00200",-- 32
x"ff800",-- -128
x"ff100",-- -240
x"ffe00",-- -32
x"00300",-- 48
x"00d00",-- 208
x"00800",-- 128
x"fe400",-- -448
x"fed00",-- -304
x"00a00",-- 160
x"00900",-- 144
x"fff00",-- -16
x"00400",-- 64
x"ff800",-- -128
x"fe600",-- -416
x"fea00",-- -352
x"ffa00",-- -96
x"01200",-- 288
x"01600",-- 352
x"00100",-- 16
x"ff100",-- -240
x"ff400",-- -192
x"ffb00",-- -80
x"01500",-- 336
x"02300",-- 560
x"00600",-- 96
x"fee00",-- -288
x"ff100",-- -240
x"ffd00",-- -48
x"01500",-- 336
x"02300",-- 560
x"00c00",-- 192
x"feb00",-- -336
x"feb00",-- -336
x"00400",-- 64
x"00b00",-- 176
x"00a00",-- 160
x"00700",-- 112
x"00800",-- 128
x"00700",-- 112
x"00400",-- 64
x"00400",-- 64
x"00200",-- 32
x"00600",-- 96
x"00300",-- 48
x"00d00",-- 208
x"01a00",-- 416
x"00100",-- 16
x"fef00",-- -272
x"00100",-- 16
x"01b00",-- 432
x"02000",-- 512
x"00900",-- 144
x"00100",-- 16
x"01400",-- 320
x"02100",-- 528
x"02200",-- 544
x"01d00",-- 464
x"00700",-- 112
x"ff600",-- -160
x"00400",-- 64
x"01b00",-- 432
x"02a00",-- 672
x"02900",-- 656
x"00a00",-- 160
x"fe400",-- -448
x"ffb00",-- -80
x"01300",-- 304
x"01600",-- 352
x"01b00",-- 432
x"00b00",-- 176
x"00000",-- 0
x"00300",-- 48
x"ffd00",-- -48
x"ffb00",-- -80
x"00b00",-- 176
x"01300",-- 304
x"ffe00",-- -32
x"ffd00",-- -48
x"ffd00",-- -48
x"00100",-- 16
x"01500",-- 336
x"00700",-- 112
x"fea00",-- -352
x"feb00",-- -336
x"ffd00",-- -48
x"00d00",-- 208
x"01100",-- 272
x"ff300",-- -208
x"fd800",-- -640
x"fd800",-- -640
x"fd600",-- -672
x"fe100",-- -496
x"ff700",-- -144
x"feb00",-- -336
x"fd600",-- -672
x"fd400",-- -704
x"fd000",-- -768
x"fcd00",-- -816
x"fcf00",-- -784
x"fcd00",-- -816
x"fce00",-- -800
x"fdb00",-- -592
x"fd700",-- -656
x"fce00",-- -800
x"fd200",-- -736
x"fdd00",-- -560
x"fd200",-- -736
x"fcc00",-- -832
x"fdc00",-- -576
x"fe000",-- -512
x"fd900",-- -624
x"fcf00",-- -784
x"fcc00",-- -832
x"fde00",-- -544
x"fe900",-- -368
x"feb00",-- -336
x"fe600",-- -416
x"fe200",-- -480
x"fdd00",-- -560
x"fdf00",-- -528
x"ff400",-- -192
x"ff800",-- -128
x"ff800",-- -128
x"00300",-- 48
x"00000",-- 0
x"ff500",-- -176
x"ff600",-- -160
x"ff400",-- -192
x"fed00",-- -304
x"ffd00",-- -48
x"01100",-- 272
x"02000",-- 512
x"01f00",-- 496
x"01900",-- 400
x"02500",-- 592
x"02400",-- 576
x"01800",-- 384
x"02300",-- 560
x"03400",-- 832
x"03600",-- 864
x"03400",-- 832
x"02f00",-- 752
x"02800",-- 640
x"02a00",-- 672
x"03200",-- 800
x"03e00",-- 992
x"04400",-- 1088
x"03d00",-- 976
x"03700",-- 880
x"04200",-- 1056
x"04e00",-- 1248
x"05a00",-- 1440
x"05f00",-- 1520
x"04900",-- 1168
x"03900",-- 912
x"05100",-- 1296
x"07300",-- 1840
x"07500",-- 1872
x"06800",-- 1664
x"06400",-- 1600
x"05b00",-- 1456
x"04a00",-- 1184
x"05400",-- 1344
x"05800",-- 1408
x"04900",-- 1168
x"04200",-- 1056
x"05200",-- 1312
x"05f00",-- 1520
x"05500",-- 1360
x"04f00",-- 1264
x"05400",-- 1344
x"04f00",-- 1264
x"02100",-- 528
x"ff300",-- -208
x"ffd00",-- -48
x"00f00",-- 240
x"ff500",-- -176
x"fc900",-- -880
x"fbd00",-- -1072
x"fa900",-- -1392
x"f8700",-- -1936
x"f6600",-- -2464
x"f6300",-- -2512
x"f7000",-- -2304
x"f7100",-- -2288
x"f6e00",-- -2336
x"f6600",-- -2464
x"f5e00",-- -2592
x"f6e00",-- -2336
x"f7800",-- -2176
x"f5e00",-- -2592
x"f4c00",-- -2880
x"f6000",-- -2560
x"f8a00",-- -1888
x"fa800",-- -1408
x"f9800",-- -1664
x"f8100",-- -2032
x"f7f00",-- -2064
x"f8d00",-- -1840
x"fad00",-- -1328
x"fc700",-- -912
x"fc000",-- -1024
x"fa400",-- -1472
x"f9500",-- -1712
x"f9c00",-- -1600
x"fb000",-- -1280
x"fb500",-- -1200
x"fa100",-- -1520
x"f9c00",-- -1600
x"fb300",-- -1232
x"fbc00",-- -1088
x"fc300",-- -976
x"fc500",-- -944
x"fbd00",-- -1072
x"fc700",-- -912
x"fe500",-- -432
x"ff300",-- -208
x"ff200",-- -224
x"ffc00",-- -64
x"00900",-- 144
x"01c00",-- 448
x"02a00",-- 672
x"02600",-- 608
x"02700",-- 624
x"03700",-- 880
x"04c00",-- 1216
x"05e00",-- 1504
x"05c00",-- 1472
x"05300",-- 1328
x"05c00",-- 1472
x"07500",-- 1872
x"08900",-- 2192
x"08000",-- 2048
x"07000",-- 1792
x"06a00",-- 1696
x"06e00",-- 1760
x"07400",-- 1856
x"08300",-- 2096
x"08d00",-- 2256
x"07e00",-- 2016
x"08000",-- 2048
x"09d00",-- 2512
x"0ad00",-- 2768
x"0ae00",-- 2784
x"09c00",-- 2496
x"09100",-- 2320
x"0a600",-- 2656
x"0ae00",-- 2784
x"0b400",-- 2880
x"0bb00",-- 2992
x"0bc00",-- 3008
x"09a00",-- 2464
x"08700",-- 2160
x"09f00",-- 2544
x"0a300",-- 2608
x"08800",-- 2176
x"09500",-- 2384
x"09e00",-- 2528
x"07900",-- 1936
x"03c00",-- 960
x"02f00",-- 752
x"03800",-- 896
x"ffb00",-- -80
x"fcd00",-- -816
x"fa800",-- -1408
x"f9200",-- -1760
x"f8e00",-- -1824
x"f8200",-- -2016
x"f7500",-- -2224
x"f5900",-- -2672
x"f3900",-- -3184
x"f2700",-- -3472
x"f3000",-- -3328
x"f3900",-- -3184
x"f1e00",-- -3616
x"f0500",-- -4016
x"ef700",-- -4240
x"f1500",-- -3760
x"f6100",-- -2544
x"f7a00",-- -2144
x"f6600",-- -2464
x"f4900",-- -2928
x"f5000",-- -2816
x"f7800",-- -2176
x"fa300",-- -1488
x"fac00",-- -1344
x"f9400",-- -1728
x"f8c00",-- -1856
x"f8b00",-- -1872
x"f9000",-- -1792
x"f9800",-- -1664
x"f9000",-- -1792
x"f8100",-- -2032
x"f7d00",-- -2096
x"f8000",-- -2048
x"f9100",-- -1776
x"f9200",-- -1760
x"f8c00",-- -1856
x"f8d00",-- -1840
x"f9300",-- -1744
x"fa900",-- -1392
x"fc000",-- -1024
x"fc800",-- -896
x"fcb00",-- -848
x"fdc00",-- -576
x"ff100",-- -240
x"ffe00",-- -32
x"00700",-- 112
x"00f00",-- 240
x"02d00",-- 720
x"04f00",-- 1264
x"05900",-- 1424
x"05e00",-- 1504
x"06200",-- 1568
x"05f00",-- 1520
x"06700",-- 1648
x"07100",-- 1808
x"07f00",-- 2032
x"08e00",-- 2272
x"08f00",-- 2288
x"08900",-- 2192
x"08800",-- 2176
x"08f00",-- 2288
x"0a100",-- 2576
x"0bd00",-- 3024
x"0c300",-- 3120
x"0b500",-- 2896
x"0b000",-- 2816
x"0bf00",-- 3056
x"0d500",-- 3408
x"0eb00",-- 3760
x"0f300",-- 3888
x"0f400",-- 3904
x"0eb00",-- 3760
x"0e500",-- 3664
x"0f000",-- 3840
x"0dd00",-- 3536
x"0d400",-- 3392
x"0ea00",-- 3744
x"10900",-- 4240
x"12100",-- 4624
x"11200",-- 4384
x"0fc00",-- 4032
x"0d200",-- 3360
x"09600",-- 2400
x"03b00",-- 944
x"00100",-- 16
x"ff400",-- -192
x"fd200",-- -736
x"faa00",-- -1376
x"f9e00",-- -1568
x"f6a00",-- -2400
x"f1e00",-- -3616
x"f0f00",-- -3856
x"f2600",-- -3488
x"f1f00",-- -3600
x"f0500",-- -4016
x"f1a00",-- -3680
x"f3000",-- -3328
x"f3800",-- -3200
x"f4100",-- -3056
x"f3f00",-- -3088
x"f3600",-- -3232
x"f5500",-- -2736
x"f7700",-- -2192
x"f7600",-- -2208
x"f7800",-- -2176
x"f8c00",-- -1856
x"f7e00",-- -2080
x"f6900",-- -2416
x"f7700",-- -2192
x"f6b00",-- -2384
x"f5e00",-- -2592
x"f6b00",-- -2384
x"f6b00",-- -2384
x"f5500",-- -2736
x"f3e00",-- -3104
x"f3500",-- -3248
x"f3400",-- -3264
x"f4200",-- -3040
x"f6000",-- -2560
x"f6500",-- -2480
x"f6800",-- -2432
x"f7300",-- -2256
x"f8000",-- -2048
x"f9300",-- -1744
x"fa400",-- -1472
x"fbc00",-- -1088
x"fc100",-- -1008
x"fd200",-- -736
x"fdf00",-- -528
x"fe000",-- -512
x"fee00",-- -288
x"00700",-- 112
x"01400",-- 320
x"02500",-- 592
x"02f00",-- 752
x"03000",-- 768
x"03500",-- 848
x"04900",-- 1168
x"05600",-- 1376
x"06500",-- 1616
x"07400",-- 1856
x"07a00",-- 1952
x"07d00",-- 2000
x"08100",-- 2064
x"09400",-- 2368
x"0a300",-- 2608
x"0a200",-- 2592
x"0ac00",-- 2752
x"0c500",-- 3152
x"0cb00",-- 3248
x"0ce00",-- 3296
x"0d500",-- 3408
x"0eb00",-- 3760
x"0f900",-- 3984
x"10c00",-- 4288
x"11d00",-- 4560
x"11100",-- 4368
x"11900",-- 4496
x"14000",-- 5120
x"17100",-- 5904
x"16200",-- 5664
x"10400",-- 4160
x"0f900",-- 3984
x"14600",-- 5216
x"19500",-- 6480
x"16b00",-- 5808
x"0a400",-- 2624
x"fff00",-- -16
x"fb900",-- -1136
x"ff100",-- -240
x"ff700",-- -144
x"fa600",-- -1440
x"f5500",-- -2736
x"f0500",-- -4016
x"ee600",-- -4512
x"ef100",-- -4336
x"f1100",-- -3824
x"ef600",-- -4256
x"eb100",-- -5360
x"ec600",-- -5024
x"f2800",-- -3456
x"f5d00",-- -2608
x"f7b00",-- -2128
x"f6800",-- -2432
x"f7000",-- -2304
x"f9600",-- -1696
x"fce00",-- -800
x"ff100",-- -240
x"fd900",-- -624
x"fd300",-- -720
x"fca00",-- -864
x"fcd00",-- -816
x"fc100",-- -1008
x"f9d00",-- -1584
x"f7100",-- -2288
x"f4c00",-- -2880
x"f3a00",-- -3168
x"f3100",-- -3312
x"f0500",-- -4016
x"eea00",-- -4448
x"eeb00",-- -4432
x"f1800",-- -3712
x"f3e00",-- -3104
x"f4500",-- -2992
x"f5400",-- -2752
x"f4e00",-- -2848
x"f6700",-- -2448
x"f9400",-- -1728
x"fc600",-- -928
x"fdd00",-- -560
x"fe000",-- -512
x"fee00",-- -288
x"fff00",-- -16
x"00600",-- 96
x"01200",-- 288
x"00d00",-- 208
x"00f00",-- 240
x"01c00",-- 448
x"02800",-- 640
x"03100",-- 784
x"02500",-- 592
x"02100",-- 528
x"02000",-- 512
x"03300",-- 816
x"04700",-- 1136
x"05000",-- 1280
x"04f00",-- 1264
x"05500",-- 1360
x"06d00",-- 1744
x"08d00",-- 2256
x"0a100",-- 2576
x"0b600",-- 2912
x"0c800",-- 3200
x"0d500",-- 3408
x"0e900",-- 3728
x"0f000",-- 3840
x"0fc00",-- 4032
x"10100",-- 4112
x"11000",-- 4352
x"11400",-- 4416
x"12100",-- 4624
x"13a00",-- 5024
x"16400",-- 5696
x"18400",-- 6208
x"19400",-- 6464
x"17f00",-- 6128
x"16a00",-- 5792
x"16b00",-- 5808
x"16000",-- 5632
x"0fe00",-- 4064
x"04b00",-- 1200
x"fc100",-- -1008
x"fa600",-- -1440
x"fc900",-- -880
x"faf00",-- -1296
x"f5c00",-- -2624
x"edc00",-- -4672
x"ea100",-- -5616
x"e9400",-- -5824
x"eb600",-- -5280
x"ec500",-- -5040
x"eb200",-- -5344
x"ecf00",-- -4880
x"f0500",-- -4016
x"f6300",-- -2512
x"fa700",-- -1424
x"fba00",-- -1120
x"fbd00",-- -1072
x"fd300",-- -720
x"00c00",-- 192
x"04d00",-- 1232
x"05a00",-- 1440
x"05500",-- 1360
x"02d00",-- 720
x"00d00",-- 208
x"feb00",-- -336
x"fc200",-- -992
x"f9700",-- -1680
x"f5800",-- -2688
x"f3300",-- -3280
x"f1300",-- -3792
x"ef500",-- -4272
x"ed600",-- -4768
x"eca00",-- -4960
x"edd00",-- -4656
x"f0600",-- -4000
x"f3100",-- -3312
x"f5100",-- -2800
x"f6000",-- -2560
x"f7b00",-- -2128
x"f9b00",-- -1616
x"fb700",-- -1168
x"fc000",-- -1024
x"fd100",-- -752
x"ffa00",-- -96
x"02200",-- 544
x"02b00",-- 688
x"01500",-- 336
x"00100",-- 16
x"ffa00",-- -96
x"00d00",-- 208
x"01f00",-- 496
x"01f00",-- 496
x"00600",-- 96
x"ff100",-- -240
x"ff400",-- -192
x"00700",-- 112
x"01800",-- 384
x"01c00",-- 448
x"01700",-- 368
x"01f00",-- 496
x"03800",-- 896
x"05200",-- 1312
x"06b00",-- 1712
x"07800",-- 1920
x"08f00",-- 2288
x"0a900",-- 2704
x"0d600",-- 3424
x"0eb00",-- 3760
x"0f200",-- 3872
x"0f600",-- 3936
x"10600",-- 4192
x"11200",-- 4384
x"10f00",-- 4336
x"11e00",-- 4576
x"11e00",-- 4576
x"14100",-- 5136
x"16100",-- 5648
x"19000",-- 6400
x"19000",-- 6400
x"18900",-- 6288
x"1aa00",-- 6816
x"1b200",-- 6944
x"15800",-- 5504
x"07c00",-- 1984
x"f7f00",-- -2064
x"f2500",-- -3504
x"f4900",-- -2928
x"f8300",-- -2000
x"f7300",-- -2256
x"f1800",-- -3712
x"ebd00",-- -5168
x"e4800",-- -7040
x"e4800",-- -7040
x"e8500",-- -6064
x"eb100",-- -5360
x"ec500",-- -5040
x"ef600",-- -4256
x"f6200",-- -2528
x"fb000",-- -1280
x"fd600",-- -672
x"feb00",-- -336
x"ff700",-- -144
x"02200",-- 544
x"07300",-- 1840
x"0b500",-- 2896
x"0c200",-- 3104
x"07900",-- 1936
x"04200",-- 1056
x"01e00",-- 480
x"00d00",-- 208
x"fd200",-- -736
x"f7e00",-- -2080
x"f4000",-- -3072
x"f0c00",-- -3904
x"ee700",-- -4496
x"ec400",-- -5056
x"eb000",-- -5376
x"eb900",-- -5232
x"ed400",-- -4800
x"f0e00",-- -3872
x"f4300",-- -3024
x"f6500",-- -2480
x"f6000",-- -2560
x"f5b00",-- -2640
x"fa900",-- -1392
x"00b00",-- 176
x"04b00",-- 1200
x"04000",-- 1024
x"02400",-- 576
x"00200",-- 32
x"fea00",-- -352
x"00600",-- 96
x"01a00",-- 416
x"02000",-- 512
x"01500",-- 336
x"00900",-- 144
x"ff900",-- -112
x"fe200",-- -480
x"fd500",-- -688
x"fc900",-- -880
x"fca00",-- -864
x"fe600",-- -416
x"ffc00",-- -64
x"00b00",-- 176
x"00800",-- 128
x"00f00",-- 240
x"02200",-- 544
x"03c00",-- 960
x"06100",-- 1552
x"07700",-- 1904
x"09700",-- 2416
x"0a900",-- 2704
x"0b600",-- 2912
x"0bb00",-- 2992
x"0c400",-- 3136
x"0df00",-- 3568
x"0ff00",-- 4080
x"11100",-- 4368
x"10500",-- 4176
x"0e800",-- 3712
x"0e200",-- 3616
x"0fe00",-- 4064
x"13200",-- 4896
x"15c00",-- 5568
x"16900",-- 5776
x"17b00",-- 6064
x"19200",-- 6432
x"1bd00",-- 7120
x"1a600",-- 6752
x"11000",-- 4352
x"fee00",-- -288
x"f0900",-- -3952
x"ef900",-- -4208
x"f5100",-- -2800
x"f7700",-- -2192
x"f4000",-- -3072
x"f0500",-- -4016
x"ec400",-- -5056
x"e8b00",-- -5968
x"e9400",-- -5824
x"eb800",-- -5248
x"eeb00",-- -4432
x"f3900",-- -3184
x"f9e00",-- -1568
x"00700",-- 112
x"03200",-- 800
x"03000",-- 768
x"01f00",-- 496
x"02900",-- 656
x"06d00",-- 1744
x"0a500",-- 2640
x"0a300",-- 2608
x"06500",-- 1616
x"03000",-- 768
x"00e00",-- 224
x"fc300",-- -976
x"f5100",-- -2800
x"f0300",-- -4048
x"eeb00",-- -4432
x"ee200",-- -4576
x"eb800",-- -5248
x"ea400",-- -5568
x"ea500",-- -5552
x"eaf00",-- -5392
x"ee800",-- -4480
x"f3b00",-- -3152
x"f8b00",-- -1872
x"fb300",-- -1232
x"fd200",-- -736
x"ff600",-- -160
x"01000",-- 256
x"02d00",-- 720
x"03b00",-- 944
x"03a00",-- 928
x"02400",-- 576
x"01300",-- 304
x"01700",-- 368
x"00d00",-- 208
x"ff700",-- -144
x"fc700",-- -912
x"fb900",-- -1136
x"faf00",-- -1296
x"f9200",-- -1760
x"f8a00",-- -1888
x"f8a00",-- -1888
x"fad00",-- -1328
x"fc700",-- -912
x"fe200",-- -480
x"00000",-- 0
x"01200",-- 288
x"03600",-- 864
x"05000",-- 1280
x"06a00",-- 1696
x"08000",-- 2048
x"07e00",-- 2016
x"08300",-- 2096
x"08500",-- 2128
x"08c00",-- 2240
x"08300",-- 2096
x"06b00",-- 1712
x"06200",-- 1568
x"05c00",-- 1472
x"07000",-- 1792
x"07a00",-- 1952
x"07c00",-- 1984
x"08800",-- 2176
x"0a600",-- 2656
x"0cc00",-- 3264
x"0e600",-- 3680
x"0f700",-- 3952
x"11500",-- 4432
x"14500",-- 5200
x"18800",-- 6272
x"1cb00",-- 7344
x"1ed00",-- 7888
x"1e700",-- 7792
x"1cb00",-- 7344
x"18800",-- 6272
x"0bf00",-- 3056
x"fa400",-- -1472
x"ee900",-- -4464
x"ef100",-- -4336
x"f4500",-- -2992
x"f4500",-- -2992
x"f0200",-- -4064
x"eb500",-- -5296
x"e6400",-- -6592
x"e4b00",-- -6992
x"e7100",-- -6384
x"ecb00",-- -4944
x"f2700",-- -3472
x"f7200",-- -2272
x"fec00",-- -320
x"04d00",-- 1232
x"07e00",-- 2016
x"07500",-- 1872
x"06900",-- 1680
x"08900",-- 2192
x"0c000",-- 3072
x"0ef00",-- 3824
x"0e700",-- 3696
x"0a100",-- 2576
x"03500",-- 848
x"fbf00",-- -1040
x"f6900",-- -2416
x"f2200",-- -3552
x"ebe00",-- -5152
x"e6b00",-- -6480
x"e5800",-- -6784
x"e7c00",-- -6208
x"e8200",-- -6112
x"e7d00",-- -6192
x"e9a00",-- -5728
x"ed800",-- -4736
x"f3200",-- -3296
x"f9500",-- -1712
x"fe900",-- -368
x"00e00",-- 224
x"02400",-- 576
x"05100",-- 1296
x"07500",-- 1872
x"08a00",-- 2208
x"08100",-- 2064
x"06100",-- 1552
x"03000",-- 768
x"ffa00",-- -96
x"ff700",-- -144
x"fef00",-- -272
x"fe700",-- -400
x"fae00",-- -1312
x"f6d00",-- -2352
x"f5800",-- -2688
x"f6000",-- -2560
x"f9000",-- -1792
x"fa600",-- -1440
x"fac00",-- -1344
x"fb200",-- -1248
x"fd800",-- -640
x"01f00",-- 496
x"05400",-- 1344
x"06c00",-- 1728
x"07100",-- 1808
x"06a00",-- 1696
x"07900",-- 1936
x"08b00",-- 2224
x"09a00",-- 2464
x"09500",-- 2384
x"08600",-- 2144
x"08400",-- 2112
x"07800",-- 1920
x"08100",-- 2064
x"08000",-- 2048
x"08400",-- 2112
x"09500",-- 2384
x"0c200",-- 3104
x"0ea00",-- 3744
x"0fc00",-- 4032
x"0f300",-- 3888
x"0eb00",-- 3760
x"10b00",-- 4272
x"13e00",-- 5088
x"19800",-- 6528
x"1cf00",-- 7408
x"1f200",-- 7968
x"1ee00",-- 7904
x"19000",-- 6400
x"0b800",-- 2944
x"f8600",-- -1952
x"ec100",-- -5104
x"ebc00",-- -5184
x"f2900",-- -3440
x"f6900",-- -2416
x"f4f00",-- -2832
x"efb00",-- -4176
x"e8b00",-- -5968
x"e5300",-- -6864
x"e8600",-- -6048
x"ee400",-- -4544
x"f4000",-- -3072
x"fae00",-- -1312
x"03600",-- 864
x"09300",-- 2352
x"09800",-- 2432
x"08200",-- 2080
x"06400",-- 1600
x"06700",-- 1648
x"09600",-- 2400
x"0cc00",-- 3264
x"0d600",-- 3424
x"09100",-- 2320
x"03400",-- 832
x"fc600",-- -928
x"f4800",-- -2944
x"ede00",-- -4640
x"ea800",-- -5504
x"eae00",-- -5408
x"e7e00",-- -6176
x"e3f00",-- -7184
x"e4900",-- -7024
x"e8900",-- -6000
x"ed000",-- -4864
x"f0200",-- -4064
x"f5c00",-- -2624
x"fae00",-- -1312
x"fea00",-- -352
x"03900",-- 912
x"06500",-- 1616
x"06600",-- 1632
x"06000",-- 1536
x"06f00",-- 1776
x"07d00",-- 2000
x"06900",-- 1680
x"04700",-- 1136
x"00700",-- 112
x"fb800",-- -1152
x"f8200",-- -2016
x"f8200",-- -2016
x"f8d00",-- -1840
x"f9600",-- -1696
x"f9000",-- -1792
x"f6f00",-- -2320
x"f6a00",-- -2400
x"f7500",-- -2224
x"fa200",-- -1504
x"fd300",-- -720
x"fff00",-- -16
x"02a00",-- 672
x"05100",-- 1296
x"07000",-- 1792
x"07f00",-- 2032
x"07900",-- 1936
x"07900",-- 1936
x"07e00",-- 2016
x"08b00",-- 2224
x"09400",-- 2368
x"08b00",-- 2224
x"07b00",-- 1968
x"06200",-- 1568
x"05d00",-- 1488
x"06700",-- 1648
x"07700",-- 1904
x"07800",-- 1920
x"08800",-- 2176
x"0b400",-- 2880
x"0dc00",-- 3520
x"0fa00",-- 4000
x"10100",-- 4112
x"0ff00",-- 4080
x"11800",-- 4480
x"15f00",-- 5616
x"1c800",-- 7296
x"1fa00",-- 8096
x"20700",-- 8304
x"1d600",-- 7520
x"12000",-- 4608
x"feb00",-- -336
x"ee000",-- -4608
x"eb700",-- -5264
x"f0100",-- -4080
x"f4000",-- -3072
x"f5200",-- -2784
x"f3000",-- -3328
x"ed100",-- -4848
x"e7000",-- -6400
x"e8500",-- -6064
x"ee000",-- -4608
x"f2c00",-- -3392
x"f9a00",-- -1632
x"02600",-- 608
x"09300",-- 2352
x"0a200",-- 2592
x"09500",-- 2384
x"08500",-- 2128
x"05d00",-- 1488
x"06400",-- 1600
x"09400",-- 2368
x"0b700",-- 2928
x"09200",-- 2336
x"04000",-- 1024
x"fdf00",-- -528
x"f6500",-- -2480
x"eeb00",-- -4432
x"e9f00",-- -5648
x"e8b00",-- -5968
x"e9b00",-- -5712
x"e9500",-- -5808
x"e7e00",-- -6176
x"e6c00",-- -6464
x"ea300",-- -5584
x"f1600",-- -3744
x"f8000",-- -2048
x"fcd00",-- -816
x"ff300",-- -208
x"02000",-- 512
x"03f00",-- 1008
x"05f00",-- 1520
x"06900",-- 1680
x"05a00",-- 1440
x"04900",-- 1168
x"03c00",-- 960
x"02f00",-- 752
x"00900",-- 144
x"fcf00",-- -784
x"f9900",-- -1648
x"f6b00",-- -2384
x"f5f00",-- -2576
x"f7600",-- -2208
x"f9600",-- -1696
x"fa700",-- -1424
x"f9200",-- -1760
x"f8e00",-- -1824
x"f9100",-- -1776
x"fbb00",-- -1104
x"ff100",-- -240
x"03b00",-- 944
x"06700",-- 1648
x"08f00",-- 2288
x"0a400",-- 2624
x"05000",-- 1280
x"05b00",-- 1456
x"07f00",-- 2032
x"07900",-- 1936
x"07e00",-- 2016
x"05d00",-- 1488
x"05500",-- 1360
x"06000",-- 1536
x"05400",-- 1344
x"04e00",-- 1248
x"05c00",-- 1472
x"06500",-- 1616
x"06000",-- 1536
x"08a00",-- 2208
x"0cb00",-- 3248
x"0eb00",-- 3760
x"10000",-- 4096
x"10f00",-- 4336
x"11f00",-- 4592
x"14e00",-- 5344
x"19200",-- 6432
x"1d600",-- 7520
x"1ec00",-- 7872
x"1fe00",-- 8160
x"1bd00",-- 7120
x"0d600",-- 3424
x"f8c00",-- -1856
x"e9d00",-- -5680
x"e7c00",-- -6208
x"ec400",-- -5056
x"f3500",-- -3248
x"f5500",-- -2736
x"f1000",-- -3840
x"ece00",-- -4896
x"e8700",-- -6032
x"ecc00",-- -4928
x"f1a00",-- -3680
x"f4600",-- -2976
x"fe700",-- -400
x"08100",-- 2064
x"0d400",-- 3392
x"0b900",-- 2960
x"0cc00",-- 3264
x"08500",-- 2128
x"05b00",-- 1456
x"03700",-- 880
x"05f00",-- 1520
x"09d00",-- 2512
x"07300",-- 1840
x"ff500",-- -176
x"f9700",-- -1680
x"f3d00",-- -3120
x"e7900",-- -6256
x"e8600",-- -6048
x"e6900",-- -6512
x"ea400",-- -5568
x"ebb00",-- -5200
x"eb100",-- -5360
x"eb900",-- -5232
x"ec500",-- -5040
x"f4a00",-- -2912
x"fc600",-- -928
x"01500",-- 336
x"01900",-- 400
x"04100",-- 1040
x"06b00",-- 1712
x"06400",-- 1600
x"04a00",-- 1184
x"03400",-- 832
x"02000",-- 512
x"00c00",-- 192
x"ff000",-- -256
x"feb00",-- -336
x"fb800",-- -1152
x"f7700",-- -2192
x"f4e00",-- -2848
x"f5b00",-- -2640
x"f8400",-- -1984
x"f8a00",-- -1888
x"fa700",-- -1424
x"fa600",-- -1440
x"fb800",-- -1152
x"fd000",-- -768
x"ff600",-- -160
x"01d00",-- 464
x"03900",-- 912
x"07500",-- 1872
x"09100",-- 2320
x"09600",-- 2400
x"07800",-- 1920
x"05b00",-- 1456
x"05000",-- 1280
x"04900",-- 1168
x"05400",-- 1344
x"03500",-- 848
x"07c00",-- 1984
x"05f00",-- 1520
x"01d00",-- 464
x"03200",-- 800
x"03900",-- 912
x"07900",-- 1936
x"08a00",-- 2208
x"09100",-- 2320
x"0e500",-- 3664
x"10b00",-- 4272
x"10e00",-- 4320
x"12000",-- 4608
x"13900",-- 5008
x"17200",-- 5920
x"18e00",-- 6368
x"1c800",-- 7296
x"1ef00",-- 7920
x"1f100",-- 7952
x"18800",-- 6272
x"05300",-- 1328
x"efd00",-- -4144
x"e5c00",-- -6720
x"e8700",-- -6032
x"edd00",-- -4656
x"f1000",-- -3840
x"f3a00",-- -3168
x"f3300",-- -3280
x"eea00",-- -4448
x"ed300",-- -4816
x"ef500",-- -4272
x"f4400",-- -3008
x"f7600",-- -2208
x"01000",-- 256
x"0dd00",-- 3536
x"11200",-- 4384
x"10000",-- 4096
x"0b600",-- 2912
x"07400",-- 1856
x"03600",-- 864
x"01200",-- 288
x"03500",-- 848
x"04200",-- 1056
x"01200",-- 288
x"fbd00",-- -1072
x"f5f00",-- -2576
x"ef700",-- -4240
x"e7400",-- -6336
x"e4c00",-- -6976
x"e7900",-- -6256
x"ebc00",-- -5184
x"eda00",-- -4704
x"ee500",-- -4528
x"f0c00",-- -3904
x"f5000",-- -2816
x"fa800",-- -1408
x"fe600",-- -416
x"00a00",-- 160
x"03000",-- 768
x"05800",-- 1408
x"06700",-- 1648
x"05b00",-- 1456
x"03d00",-- 976
x"00700",-- 112
x"fd500",-- -688
x"fc900",-- -880
x"fd300",-- -720
x"fc500",-- -944
x"f9500",-- -1712
x"f6300",-- -2512
x"f5c00",-- -2624
x"f7600",-- -2208
x"f8700",-- -1936
x"f9a00",-- -1632
x"fb200",-- -1248
x"fc900",-- -880
x"fdf00",-- -528
x"ffa00",-- -96
x"01000",-- 256
x"02600",-- 608
x"04d00",-- 1232
x"07300",-- 1840
x"08b00",-- 2224
x"09700",-- 2416
x"08100",-- 2064
x"05700",-- 1392
x"03900",-- 912
x"03100",-- 784
x"03900",-- 912
x"03c00",-- 960
x"03a00",-- 928
x"03a00",-- 928
x"03500",-- 848
x"03f00",-- 1008
x"06400",-- 1600
x"07600",-- 1888
x"08300",-- 2096
x"0ac00",-- 2752
x"0ec00",-- 3776
x"12300",-- 4656
x"13c00",-- 5056
x"14600",-- 5216
x"14a00",-- 5280
x"15100",-- 5392
x"17f00",-- 6128
x"1c100",-- 7184
x"1d600",-- 7520
x"1c500",-- 7248
x"14000",-- 5120
x"02400",-- 576
x"ee300",-- -4560
x"e3800",-- -7296
x"e6700",-- -6544
x"eb600",-- -5280
x"eef00",-- -4368
x"f3200",-- -3296
x"f6000",-- -2560
x"f4d00",-- -2864
x"f3500",-- -3248
x"f5500",-- -2736
x"f7b00",-- -2128
x"fb700",-- -1168
x"03300",-- 816
x"0c800",-- 3200
x"11e00",-- 4576
x"10f00",-- 4336
x"0b800",-- 2944
x"05400",-- 1344
x"ff400",-- -192
x"fc600",-- -928
x"fbf00",-- -1040
x"fd100",-- -752
x"fcd00",-- -816
x"fae00",-- -1312
x"f6000",-- -2560
x"ede00",-- -4640
x"e7000",-- -6400
x"e5300",-- -6864
x"e9600",-- -5792
x"ed100",-- -4848
x"f0200",-- -4064
x"f3500",-- -3248
x"f7d00",-- -2096
x"fbf00",-- -1040
x"fe100",-- -496
x"ff500",-- -176
x"00500",-- 80
x"02000",-- 512
x"04a00",-- 1184
x"06400",-- 1600
x"05f00",-- 1520
x"01f00",-- 496
x"fd500",-- -688
x"fa100",-- -1520
x"f9000",-- -1792
x"f9b00",-- -1616
x"f8e00",-- -1824
x"f8f00",-- -1808
x"f8800",-- -1920
x"f8300",-- -2000
x"f9300",-- -1744
x"fa700",-- -1424
x"fa100",-- -1520
x"fad00",-- -1328
x"fd500",-- -688
x"00000",-- 0
x"02a00",-- 672
x"03e00",-- 992
x"05900",-- 1424
x"06900",-- 1680
x"07100",-- 1808
x"07800",-- 1920
x"07400",-- 1856
x"05b00",-- 1456
x"04200",-- 1056
x"02e00",-- 736
x"02400",-- 576
x"01600",-- 352
x"00e00",-- 224
x"01700",-- 368
x"02600",-- 608
x"04100",-- 1040
x"05200",-- 1312
x"06d00",-- 1744
x"07e00",-- 2016
x"09700",-- 2416
x"0b500",-- 2896
x"0e300",-- 3632
x"11c00",-- 4544
x"13500",-- 4944
x"14300",-- 5168
x"14900",-- 5264
x"15b00",-- 5552
x"18a00",-- 6304
x"1b700",-- 7024
x"1b800",-- 7040
x"19800",-- 6528
x"12900",-- 4752
x"05400",-- 1344
x"f2000",-- -3584
x"e5600",-- -6816
x"e5e00",-- -6688
x"e9e00",-- -5664
x"ece00",-- -4896
x"f0c00",-- -3904
x"f7500",-- -2224
x"fb300",-- -1232
x"fa300",-- -1488
x"f9d00",-- -1584
x"faa00",-- -1376
x"fba00",-- -1120
x"00600",-- 96
x"08d00",-- 2256
x"10600",-- 4192
x"10f00",-- 4336
x"0b800",-- 2944
x"05500",-- 1360
x"fe900",-- -368
x"f9500",-- -1712
x"f6a00",-- -2400
x"f7500",-- -2224
x"f8b00",-- -1872
x"f8a00",-- -1888
x"f7c00",-- -2112
x"f3c00",-- -3136
x"ee400",-- -4544
x"ea400",-- -5568
x"e9f00",-- -5648
x"ebf00",-- -5136
x"ef400",-- -4288
x"f4700",-- -2960
x"fa700",-- -1424
x"ff000",-- -256
x"00600",-- 96
x"ffb00",-- -80
x"feb00",-- -336
x"fed00",-- -304
x"00400",-- 64
x"01f00",-- 496
x"03200",-- 800
x"02700",-- 624
x"ffb00",-- -80
x"fc900",-- -880
x"f9500",-- -1712
x"f7800",-- -2176
x"f6c00",-- -2368
x"f7500",-- -2224
x"f9000",-- -1792
x"fb000",-- -1280
x"fc700",-- -912
x"fd100",-- -752
x"fc000",-- -1024
x"fa900",-- -1392
x"fba00",-- -1120
x"fe100",-- -496
x"01700",-- 368
x"04100",-- 1040
x"06800",-- 1664
x"08100",-- 2064
x"08100",-- 2064
x"06c00",-- 1728
x"04b00",-- 1200
x"03200",-- 800
x"02500",-- 592
x"02200",-- 544
x"02800",-- 640
x"02700",-- 624
x"01c00",-- 448
x"01800",-- 384
x"01100",-- 272
x"02100",-- 528
x"03700",-- 880
x"05600",-- 1376
x"08a00",-- 2208
x"0b100",-- 2832
x"0d100",-- 3344
x"0ed00",-- 3792
x"10a00",-- 4256
x"11700",-- 4464
x"12700",-- 4720
x"13200",-- 4896
x"13e00"-- 5088

);
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: top PORT MAP (
          clk => clk,
          rstn => rstn,
          i_volume => i_volume,
          i_SDATA_IN => i_SDATA_IN,
          o_SDATA_out => o_SDATA_out,
          o_SYNC => o_SYNC,
          o_RSTN => o_RSTN,
          i_BIT_CLK => i_BIT_CLK
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 
   i_BIT_CLK_process :process
   begin
		i_BIT_CLK <= '0';
		wait for i_BIT_CLK_period/2;
		i_BIT_CLK <= '1';
		wait for i_BIT_CLK_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin	
		rstn <= '0';
		-- hold reset state for 100 ns.
		wait for 100 ns;	
		rstn <= '1';
		i_volume <= (others => '1');

	wait for i_bit_clk_period*55;
		
		for j in 42 to len-1 loop
			--for k in 0 to 1 loop
				for i in 19 downto 0 loop
					i_sdata_in <= s(j)(i);
					wait for i_bit_clk_period;
				end loop;
				for i in 19 downto 0 loop
					i_sdata_in <= s(j)(i);
					wait for i_bit_clk_period;
				end loop;
			--end loop;
			wait for i_bit_clk_period*216;
		end loop;

		wait;
   end process;

END;
