--------------------------------------------------------------------------------
-- Company: 
-- Engineer: Niklas Aldn
--
-- Create Date:   17:00:43 03/25/2015
-- Design Name:   
-- Module Name:   D:/Google Drive/Exjobb/vhdl/agc_and_ac97/tb_top.vhd
-- Project Name:  agc_and_ac97
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: top
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
 
ENTITY tb_top IS
END tb_top;
 
ARCHITECTURE behavior OF tb_top IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT top
    PORT(
         clk : IN  std_logic;
         rstn : IN  std_logic;
         i_volume : IN  std_logic_vector(4 downto 0);
			i_agc_enable		: in std_logic;
         i_SDATA_IN : IN  std_logic;
         o_SDATA_out : OUT  std_logic;
         o_SYNC : OUT  std_logic;
         o_RSTN : OUT  std_logic;
         i_BIT_CLK : IN  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal rstn : std_logic := '0';
   signal i_volume : std_logic_vector(4 downto 0) := (others => '0');
	signal i_agc_enable		: std_logic := '1';
   signal i_SDATA_IN : std_logic := '0';
   signal i_BIT_CLK : std_logic := '0';

 	--Outputs
   signal o_SDATA_out : std_logic;
   signal o_SYNC : std_logic;
   signal o_RSTN : std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns; -- 100MHz
   constant i_BIT_CLK_period : time := 81.38 ns; -- 12.288 MHz
   
   constant len : integer range 0 to 65535 := 44999;
   
	type t_sample is array(19 downto 0) of std_logic;
	type t_sample_matrix is array(0 to len-1) of t_sample;
	
	signal s : t_sample_matrix := (	
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00020",-- 2
x"00020",-- 2
x"00020",-- 2
x"00000",-- 0
x"00000",-- 0
x"00020",-- 2
x"00030",-- 3
x"00030",-- 3
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00020",-- 2
x"00050",-- 5
x"00020",-- 2
x"fffe0",-- -2
x"fff80",-- -8
x"fff60",-- -10
x"fffe0",-- -2
x"00020",-- 2
x"00030",-- 3
x"00030",-- 3
x"00000",-- 0
x"fff90",-- -7
x"fff90",-- -7
x"fffd0",-- -3
x"00030",-- 3
x"000a0",-- 10
x"fffe0",-- -2
x"fff10",-- -15
x"fff90",-- -7
x"000c0",-- 12
x"000d0",-- 13
x"fff80",-- -8
x"ffdd0",-- -35
x"ffe40",-- -28
x"fffd0",-- -3
x"00070",-- 7
x"00000",-- 0
x"ffec0",-- -20
x"ffdd0",-- -35
x"ffe50",-- -27
x"00030",-- 3
x"00110",-- 17
x"00050",-- 5
x"ffee0",-- -18
x"ffea0",-- -22
x"00050",-- 5
x"00190",-- 25
x"00120",-- 18
x"00050",-- 5
x"00050",-- 5
x"000c0",-- 12
x"00170",-- 23
x"001c0",-- 28
x"001c0",-- 28
x"002b0",-- 43
x"00350",-- 53
x"00250",-- 37
x"000c0",-- 12
x"00000",-- 0
x"000f0",-- 15
x"001e0",-- 30
x"000c0",-- 12
x"fff90",-- -7
x"00020",-- 2
x"001b0",-- 27
x"00200",-- 32
x"00200",-- 32
x"00120",-- 18
x"fffe0",-- -2
x"00000",-- 0
x"00120",-- 18
x"00170",-- 23
x"000f0",-- 15
x"00000",-- 0
x"00070",-- 7
x"00160",-- 22
x"000d0",-- 13
x"00000",-- 0
x"fff90",-- -7
x"00050",-- 5
x"00170",-- 23
x"002b0",-- 43
x"00370",-- 55
x"00260",-- 38
x"000f0",-- 15
x"00000",-- 0
x"fff60",-- -10
x"fff80",-- -8
x"fff90",-- -7
x"fffe0",-- -2
x"fffd0",-- -3
x"fff80",-- -8
x"ffef0",-- -17
x"fff30",-- -13
x"00000",-- 0
x"00000",-- 0
x"fff90",-- -7
x"00000",-- 0
x"fff90",-- -7
x"fffd0",-- -3
x"002b0",-- 43
x"003e0",-- 62
x"002a0",-- 42
x"00070",-- 7
x"00080",-- 8
x"000a0",-- 10
x"001c0",-- 28
x"002b0",-- 43
x"00190",-- 25
x"00000",-- 0
x"ffec0",-- -20
x"00000",-- 0
x"000d0",-- 13
x"00000",-- 0
x"ffce0",-- -50
x"ff9c0",-- -100
x"ffae0",-- -82
x"00030",-- 3
x"003f0",-- 63
x"00210",-- 33
x"ffce0",-- -50
x"ffc10",-- -63
x"ffec0",-- -20
x"00260",-- 38
x"004b0",-- 75
x"000f0",-- 15
x"fff30",-- -13
x"ffe90",-- -23
x"000d0",-- 13
x"00370",-- 55
x"00350",-- 53
x"00000",-- 0
x"ffd30",-- -45
x"ffda0",-- -38
x"ffdf0",-- -33
x"fffe0",-- -2
x"000a0",-- 10
x"ffe00",-- -32
x"ffc40",-- -60
x"ffdf0",-- -33
x"ffd50",-- -43
x"ffec0",-- -20
x"fffb0",-- -5
x"fff60",-- -10
x"ffda0",-- -38
x"ffc70",-- -57
x"00030",-- 3
x"003e0",-- 62
x"00390",-- 57
x"fff80",-- -8
x"ffb00",-- -80
x"ffab0",-- -85
x"ffd50",-- -43
x"ffe50",-- -27
x"ffce0",-- -50
x"ff7e0",-- -130
x"ff740",-- -140
x"ffdb0",-- -37
x"003a0",-- 58
x"002f0",-- 47
x"ffc90",-- -55
x"ffa30",-- -93
x"ffdf0",-- -33
x"00300",-- 48
x"00280",-- 40
x"fff40",-- -12
x"ffe20",-- -30
x"fff40",-- -12
x"001e0",-- 30
x"002f0",-- 47
x"00120",-- 18
x"ffe90",-- -23
x"00000",-- 0
x"005f0",-- 95
x"009e0",-- 158
x"00610",-- 97
x"fff90",-- -7
x"ffbd0",-- -67
x"ffd00",-- -48
x"00080",-- 8
x"00070",-- 7
x"ffd80",-- -40
x"ffce0",-- -50
x"ffdb0",-- -37
x"ffd30",-- -45
x"ffb80",-- -72
x"ffbf0",-- -65
x"fff40",-- -12
x"000d0",-- 13
x"fffb0",-- -5
x"ffd10",-- -47
x"ffe20",-- -30
x"00000",-- 0
x"ffec0",-- -20
x"fff30",-- -13
x"00280",-- 40
x"002a0",-- 42
x"ffdb0",-- -37
x"ffb80",-- -72
x"fffd0",-- -3
x"00410",-- 65
x"00080",-- 8
x"ffdb0",-- -37
x"fff90",-- -7
x"000d0",-- 13
x"fffe0",-- -2
x"ffa10",-- -95
x"ff8b0",-- -117
x"ffea0",-- -22
x"00280",-- 40
x"00110",-- 17
x"ffd60",-- -42
x"ffd80",-- -40
x"00070",-- 7
x"00190",-- 25
x"fff80",-- -8
x"ffd00",-- -48
x"ffbd0",-- -67
x"ffe70",-- -25
x"001e0",-- 30
x"001b0",-- 27
x"ffe50",-- -27
x"ffd10",-- -47
x"ffea0",-- -22
x"fff10",-- -15
x"ffe20",-- -30
x"ffb30",-- -77
x"ff7c0",-- -132
x"ff6c0",-- -148
x"ffa60",-- -90
x"ffb50",-- -75
x"ff920",-- -110
x"ffb50",-- -75
x"ffe90",-- -23
x"ffd00",-- -48
x"ffb30",-- -77
x"ffd50",-- -43
x"fff80",-- -8
x"ffe90",-- -23
x"ffcc0",-- -52
x"ffd80",-- -40
x"00080",-- 8
x"005a0",-- 90
x"00800",-- 128
x"00530",-- 83
x"00030",-- 3
x"ffec0",-- -20
x"00140",-- 20
x"002f0",-- 47
x"00000",-- 0
x"ffc40",-- -60
x"ffc20",-- -62
x"fffe0",-- -2
x"00370",-- 55
x"00210",-- 33
x"ffd80",-- -40
x"ffa30",-- -93
x"ff990",-- -103
x"ffe00",-- -32
x"00370",-- 55
x"003e0",-- 62
x"001e0",-- 30
x"00030",-- 3
x"ffdb0",-- -37
x"ffea0",-- -22
x"00120",-- 18
x"00160",-- 22
x"001b0",-- 27
x"00210",-- 33
x"00080",-- 8
x"fffd0",-- -3
x"00000",-- 0
x"002a0",-- 42
x"00350",-- 53
x"00050",-- 5
x"ffdf0",-- -33
x"ffcb0",-- -53
x"ffd50",-- -43
x"fff40",-- -12
x"00080",-- 8
x"ffee0",-- -18
x"ffe20",-- -30
x"ffd80",-- -40
x"ffec0",-- -20
x"000c0",-- 12
x"000a0",-- 10
x"ffd50",-- -43
x"ffab0",-- -85
x"fff10",-- -15
x"00640",-- 100
x"007a0",-- 122
x"00050",-- 5
x"ff9c0",-- -100
x"ffa30",-- -93
x"ffdd0",-- -35
x"ffdd0",-- -35
x"ffb20",-- -78
x"ff9c0",-- -100
x"ffd30",-- -45
x"00000",-- 0
x"00140",-- 20
x"00070",-- 7
x"00070",-- 7
x"00020",-- 2
x"ffea0",-- -22
x"00000",-- 0
x"001e0",-- 30
x"fff90",-- -7
x"ffb20",-- -78
x"ffa90",-- -87
x"fff80",-- -8
x"004b0",-- 75
x"003f0",-- 63
x"ffea0",-- -22
x"ff9e0",-- -98
x"ffa40",-- -92
x"ffdf0",-- -33
x"ffe70",-- -25
x"ffd60",-- -42
x"ffc90",-- -55
x"ffc20",-- -62
x"ffc60",-- -58
x"ffd80",-- -40
x"ffec0",-- -20
x"00070",-- 7
x"00210",-- 33
x"00350",-- 53
x"00460",-- 70
x"002d0",-- 45
x"00110",-- 17
x"00170",-- 23
x"00610",-- 97
x"007d0",-- 125
x"00500",-- 80
x"00250",-- 37
x"000f0",-- 15
x"001b0",-- 27
x"004e0",-- 78
x"00640",-- 100
x"00280",-- 40
x"ffda0",-- -38
x"ff9e0",-- -98
x"ff9f0",-- -97
x"ffd50",-- -43
x"00000",-- 0
x"00410",-- 65
x"00440",-- 68
x"fff40",-- -12
x"ffcb0",-- -53
x"ffd60",-- -42
x"00160",-- 22
x"003e0",-- 62
x"00200",-- 32
x"fff60",-- -10
x"ffec0",-- -20
x"00020",-- 2
x"00000",-- 0
x"ffd00",-- -48
x"ffd50",-- -43
x"00030",-- 3
x"00110",-- 17
x"fffb0",-- -5
x"ffd10",-- -47
x"ffd50",-- -43
x"ffef0",-- -17
x"ffea0",-- -22
x"ffec0",-- -20
x"00070",-- 7
x"00190",-- 25
x"00160",-- 22
x"ffd80",-- -40
x"ffa80",-- -88
x"ffdb0",-- -37
x"003e0",-- 62
x"00800",-- 128
x"00570",-- 87
x"001c0",-- 28
x"fffb0",-- -5
x"002f0",-- 47
x"007a0",-- 122
x"004b0",-- 75
x"fff40",-- -12
x"ffd80",-- -40
x"00210",-- 33
x"006c0",-- 108
x"00370",-- 55
x"ffd80",-- -40
x"ffea0",-- -22
x"003c0",-- 60
x"00640",-- 100
x"00570",-- 87
x"00480",-- 72
x"003e0",-- 62
x"00230",-- 35
x"00160",-- 22
x"00410",-- 65
x"00840",-- 132
x"00940",-- 148
x"004d0",-- 77
x"001b0",-- 27
x"00210",-- 33
x"00350",-- 53
x"00390",-- 57
x"00120",-- 18
x"00030",-- 3
x"00000",-- 0
x"000c0",-- 12
x"00300",-- 48
x"00210",-- 33
x"ffea0",-- -22
x"ffc20",-- -62
x"ffda0",-- -38
x"001e0",-- 30
x"00410",-- 65
x"00110",-- 17
x"ffc40",-- -60
x"ffbc0",-- -68
x"ffef0",-- -17
x"003a0",-- 58
x"00550",-- 85
x"00260",-- 38
x"000c0",-- 12
x"002b0",-- 43
x"00320",-- 50
x"fff80",-- -8
x"ffb00",-- -80
x"ffa90",-- -87
x"ffc60",-- -58
x"ffc90",-- -55
x"ffcc0",-- -52
x"ffbc0",-- -68
x"ffd80",-- -40
x"00230",-- 35
x"00430",-- 67
x"fffb0",-- -5
x"ff950",-- -107
x"ffce0",-- -50
x"00550",-- 85
x"00730",-- 115
x"00350",-- 53
x"00020",-- 2
x"00070",-- 7
x"00320",-- 50
x"005f0",-- 95
x"005f0",-- 95
x"00350",-- 53
x"00160",-- 22
x"00080",-- 8
x"00230",-- 35
x"00430",-- 67
x"00300",-- 48
x"fff40",-- -12
x"ffce0",-- -50
x"ffee0",-- -18
x"fff40",-- -12
x"ffe00",-- -32
x"ffdf0",-- -33
x"ffe20",-- -30
x"ffce0",-- -50
x"ffc90",-- -55
x"ffd80",-- -40
x"00000",-- 0
x"00390",-- 57
x"00440",-- 68
x"00080",-- 8
x"fff40",-- -12
x"00210",-- 33
x"002a0",-- 42
x"00080",-- 8
x"ffe50",-- -27
x"ffe70",-- -25
x"00000",-- 0
x"fff90",-- -7
x"ffdf0",-- -33
x"ffd30",-- -45
x"ffef0",-- -17
x"00080",-- 8
x"00080",-- 8
x"00000",-- 0
x"ffda0",-- -38
x"ffe00",-- -32
x"fff60",-- -10
x"00080",-- 8
x"00050",-- 5
x"fff40",-- -12
x"00000",-- 0
x"fff90",-- -7
x"00050",-- 5
x"fffe0",-- -2
x"ffdb0",-- -37
x"ffec0",-- -20
x"001c0",-- 28
x"001b0",-- 27
x"fff30",-- -13
x"ffd10",-- -47
x"ffcc0",-- -52
x"ffe50",-- -27
x"fff80",-- -8
x"fff30",-- -13
x"ffbc0",-- -68
x"ffdf0",-- -33
x"002d0",-- 45
x"001b0",-- 27
x"ffcb0",-- -53
x"ffc20",-- -62
x"002b0",-- 43
x"00930",-- 147
x"00660",-- 102
x"ffec0",-- -20
x"ff9c0",-- -100
x"ffd00",-- -48
x"003a0",-- 58
x"003a0",-- 58
x"ffdf0",-- -33
x"ffad0",-- -83
x"ffd50",-- -43
x"000f0",-- 15
x"00250",-- 37
x"fff60",-- -10
x"ffad0",-- -83
x"ffab0",-- -85
x"ffe50",-- -27
x"ffdd0",-- -35
x"ff900",-- -112
x"ff670",-- -153
x"ff990",-- -103
x"fff40",-- -12
x"00250",-- 37
x"00120",-- 18
x"ffee0",-- -18
x"ffea0",-- -22
x"00020",-- 2
x"002f0",-- 47
x"003e0",-- 62
x"00320",-- 50
x"001e0",-- 30
x"00000",-- 0
x"ffdf0",-- -33
x"ffec0",-- -20
x"00300",-- 48
x"003c0",-- 60
x"00020",-- 2
x"ffbc0",-- -68
x"ffb80",-- -72
x"ffef0",-- -17
x"00000",-- 0
x"00020",-- 2
x"fff10",-- -15
x"ffe00",-- -32
x"fffe0",-- -2
x"00280",-- 40
x"003a0",-- 58
x"001e0",-- 30
x"00050",-- 5
x"00110",-- 17
x"fffd0",-- -3
x"ffd60",-- -42
x"ffdf0",-- -33
x"00070",-- 7
x"00320",-- 50
x"000f0",-- 15
x"ffda0",-- -38
x"ffc20",-- -62
x"ffea0",-- -22
x"00280",-- 40
x"00480",-- 72
x"00170",-- 23
x"ffda0",-- -38
x"ffcc0",-- -52
x"ffec0",-- -20
x"003a0",-- 58
x"00370",-- 55
x"ffef0",-- -17
x"ffc70",-- -57
x"ffe40",-- -28
x"00000",-- 0
x"ffe40",-- -28
x"ffe20",-- -30
x"00000",-- 0
x"003a0",-- 58
x"004b0",-- 75
x"fffb0",-- -5
x"ffbc0",-- -68
x"ffc90",-- -55
x"ffee0",-- -18
x"fff40",-- -12
x"ffdd0",-- -35
x"ffce0",-- -50
x"ffdf0",-- -33
x"002a0",-- 42
x"00640",-- 100
x"00620",-- 98
x"004b0",-- 75
x"00120",-- 18
x"ffd80",-- -40
x"ffb80",-- -72
x"ffef0",-- -17
x"00410",-- 65
x"00530",-- 83
x"00210",-- 33
x"fffe0",-- -2
x"00000",-- 0
x"001e0",-- 30
x"00490",-- 73
x"00440",-- 68
x"001e0",-- 30
x"000f0",-- 15
x"003f0",-- 63
x"00500",-- 80
x"005d0",-- 93
x"004d0",-- 77
x"00280",-- 40
x"00350",-- 53
x"00280",-- 40
x"002a0",-- 42
x"00390",-- 57
x"002f0",-- 47
x"fff80",-- -8
x"ffd30",-- -45
x"ffe70",-- -25
x"000c0",-- 12
x"004d0",-- 77
x"00410",-- 65
x"ffea0",-- -22
x"ffa90",-- -87
x"ffa40",-- -92
x"ffdf0",-- -33
x"fffb0",-- -5
x"00020",-- 2
x"001b0",-- 27
x"00160",-- 22
x"00000",-- 0
x"ffe00",-- -32
x"fff10",-- -15
x"00170",-- 23
x"00520",-- 82
x"005d0",-- 93
x"001b0",-- 27
x"fff90",-- -7
x"00120",-- 18
x"002f0",-- 47
x"00250",-- 37
x"00080",-- 8
x"ffea0",-- -22
x"ffe90",-- -23
x"fff80",-- -8
x"00210",-- 33
x"00250",-- 37
x"fff10",-- -15
x"ffd10",-- -47
x"ffe20",-- -30
x"00230",-- 35
x"005c0",-- 92
x"00440",-- 68
x"00020",-- 2
x"fff40",-- -12
x"000a0",-- 10
x"00120",-- 18
x"00280",-- 40
x"00350",-- 53
x"00190",-- 25
x"ffd10",-- -47
x"ffc40",-- -60
x"fffd0",-- -3
x"002f0",-- 47
x"001b0",-- 27
x"00020",-- 2
x"00200",-- 32
x"00480",-- 72
x"00490",-- 73
x"fff60",-- -10
x"ffbd0",-- -67
x"ffd10",-- -47
x"001b0",-- 27
x"00370",-- 55
x"00000",-- 0
x"ffd50",-- -43
x"ffdb0",-- -37
x"ffd80",-- -40
x"ffc60",-- -58
x"ffd00",-- -48
x"ffd60",-- -42
x"ffec0",-- -20
x"ffee0",-- -18
x"ffd80",-- -40
x"ffcb0",-- -53
x"ffbc0",-- -68
x"ffcc0",-- -52
x"fff10",-- -15
x"fff30",-- -13
x"ffe40",-- -28
x"ffb70",-- -73
x"ffab0",-- -85
x"ffd60",-- -42
x"ffec0",-- -20
x"ffe20",-- -30
x"ffc70",-- -57
x"ffc10",-- -63
x"ffc90",-- -55
x"ffdf0",-- -33
x"00030",-- 3
x"fff10",-- -15
x"ffa10",-- -95
x"ffa30",-- -93
x"ffe20",-- -30
x"001e0",-- 30
x"00080",-- 8
x"ffb80",-- -72
x"ffa90",-- -87
x"ffce0",-- -50
x"fff10",-- -15
x"ffe00",-- -32
x"ffdf0",-- -33
x"ffea0",-- -22
x"fffb0",-- -5
x"fff80",-- -8
x"ffea0",-- -22
x"fff80",-- -8
x"00000",-- 0
x"fff90",-- -7
x"ffe70",-- -25
x"ffbf0",-- -65
x"ff9a0",-- -102
x"ffbd0",-- -67
x"00000",-- 0
x"00260",-- 38
x"fffd0",-- -3
x"ffb50",-- -75
x"ffab0",-- -85
x"fff60",-- -10
x"001b0",-- 27
x"00000",-- 0
x"ffc40",-- -60
x"ff920",-- -110
x"ffba0",-- -70
x"00080",-- 8
x"00170",-- 23
x"fffb0",-- -5
x"ffdf0",-- -33
x"ffc60",-- -58
x"ffbf0",-- -65
x"ffc20",-- -62
x"ffcc0",-- -52
x"ffc40",-- -60
x"ffc20",-- -62
x"ffd80",-- -40
x"ffdf0",-- -33
x"ffce0",-- -50
x"ffbc0",-- -68
x"ffe70",-- -25
x"001e0",-- 30
x"001e0",-- 30
x"00000",-- 0
x"fff40",-- -12
x"fffd0",-- -3
x"00160",-- 22
x"00260",-- 38
x"fffd0",-- -3
x"ffc60",-- -58
x"ffbc0",-- -68
x"ffec0",-- -20
x"002f0",-- 47
x"004b0",-- 75
x"00500",-- 80
x"002b0",-- 43
x"00050",-- 5
x"00080",-- 8
x"00250",-- 37
x"00570",-- 87
x"00610",-- 97
x"002f0",-- 47
x"fff40",-- -12
x"ffdf0",-- -33
x"00080",-- 8
x"005f0",-- 95
x"00610",-- 97
x"00260",-- 38
x"fffd0",-- -3
x"fff40",-- -12
x"00370",-- 55
x"00700",-- 112
x"00440",-- 68
x"fffb0",-- -5
x"ffea0",-- -22
x"00080",-- 8
x"00280",-- 40
x"000a0",-- 10
x"fff10",-- -15
x"ffdf0",-- -33
x"00020",-- 2
x"00210",-- 33
x"001e0",-- 30
x"00320",-- 50
x"003a0",-- 58
x"00140",-- 20
x"ffc10",-- -63
x"ff970",-- -105
x"ffea0",-- -22
x"003e0",-- 62
x"00300",-- 48
x"ffea0",-- -22
x"ffa30",-- -93
x"ffbc0",-- -68
x"00030",-- 3
x"002a0",-- 42
x"00210",-- 33
x"fff40",-- -12
x"ffd30",-- -45
x"fff10",-- -15
x"003a0",-- 58
x"00520",-- 82
x"00210",-- 33
x"ffe70",-- -25
x"ffda0",-- -38
x"00190",-- 25
x"005c0",-- 92
x"00490",-- 73
x"fffb0",-- -5
x"ffd80",-- -40
x"ffee0",-- -18
x"00000",-- 0
x"000a0",-- 10
x"00120",-- 18
x"00250",-- 37
x"001b0",-- 27
x"ffec0",-- -20
x"ffbf0",-- -65
x"ffea0",-- -22
x"001b0",-- 27
x"00020",-- 2
x"ffbd0",-- -67
x"ffa30",-- -93
x"ffda0",-- -38
x"fff80",-- -8
x"fff30",-- -13
x"ffdb0",-- -37
x"ffea0",-- -22
x"ffee0",-- -18
x"ffe70",-- -25
x"00020",-- 2
x"00070",-- 7
x"fffe0",-- -2
x"fff30",-- -13
x"fff80",-- -8
x"00160",-- 22
x"00440",-- 68
x"001b0",-- 27
x"ffd10",-- -47
x"ffc90",-- -55
x"fffe0",-- -2
x"001b0",-- 27
x"fff60",-- -10
x"ffb50",-- -75
x"ff800",-- -128
x"ff970",-- -105
x"ffd00",-- -48
x"fff10",-- -15
x"ffc70",-- -57
x"ff830",-- -125
x"ff860",-- -122
x"ffa90",-- -87
x"ffa80",-- -88
x"ff9f0",-- -97
x"ff7e0",-- -130
x"ff670",-- -153
x"ff800",-- -128
x"ffb80",-- -72
x"ffef0",-- -17
x"fff80",-- -8
x"00020",-- 2
x"ffef0",-- -17
x"ffd60",-- -42
x"ffdf0",-- -33
x"ffec0",-- -20
x"fff10",-- -15
x"000c0",-- 12
x"001c0",-- 28
x"ffef0",-- -17
x"ffb80",-- -72
x"ffc10",-- -63
x"00050",-- 5
x"003a0",-- 58
x"00370",-- 55
x"00050",-- 5
x"fff80",-- -8
x"001b0",-- 27
x"00480",-- 72
x"001e0",-- 30
x"ffec0",-- -20
x"fffe0",-- -2
x"00160",-- 22
x"001b0",-- 27
x"00250",-- 37
x"002b0",-- 43
x"00050",-- 5
x"ffe50",-- -27
x"ffd80",-- -40
x"00140",-- 20
x"00480",-- 72
x"001e0",-- 30
x"ffbf0",-- -65
x"ffa10",-- -95
x"ffe50",-- -27
x"00210",-- 33
x"001b0",-- 27
x"ffd10",-- -47
x"ffb70",-- -73
x"ffc60",-- -58
x"ffdf0",-- -33
x"ffea0",-- -22
x"000c0",-- 12
x"00340",-- 52
x"001b0",-- 27
x"fff10",-- -15
x"ffdf0",-- -33
x"ffe50",-- -27
x"ffee0",-- -18
x"001c0",-- 28
x"00200",-- 32
x"00170",-- 23
x"002b0",-- 43
x"00260",-- 38
x"002f0",-- 47
x"00280",-- 40
x"000c0",-- 12
x"000c0",-- 12
x"00210",-- 33
x"002f0",-- 47
x"00190",-- 25
x"ffea0",-- -22
x"ffe20",-- -30
x"00000",-- 0
x"00170",-- 23
x"00120",-- 18
x"00170",-- 23
x"00160",-- 22
x"00110",-- 17
x"00020",-- 2
x"000f0",-- 15
x"002b0",-- 43
x"00250",-- 37
x"003a0",-- 58
x"003a0",-- 58
x"003a0",-- 58
x"002f0",-- 47
x"004b0",-- 75
x"00670",-- 103
x"00780",-- 120
x"00670",-- 103
x"00280",-- 40
x"00200",-- 32
x"00340",-- 52
x"00500",-- 80
x"00320",-- 50
x"000c0",-- 12
x"00210",-- 33
x"00570",-- 87
x"00440",-- 68
x"00050",-- 5
x"fff60",-- -10
x"00080",-- 8
x"002b0",-- 43
x"002f0",-- 47
x"00110",-- 17
x"ffec0",-- -20
x"ffce0",-- -50
x"ffbf0",-- -65
x"ffc90",-- -55
x"fff60",-- -10
x"00110",-- 17
x"00030",-- 3
x"ffef0",-- -17
x"ffef0",-- -17
x"fff40",-- -12
x"00050",-- 5
x"00000",-- 0
x"ffda0",-- -38
x"ffd50",-- -43
x"ffdb0",-- -37
x"ffe20",-- -30
x"ffd80",-- -40
x"ffe40",-- -28
x"000c0",-- 12
x"00210",-- 33
x"ffea0",-- -22
x"ffdf0",-- -33
x"ffe50",-- -27
x"ffdf0",-- -33
x"fffe0",-- -2
x"000c0",-- 12
x"000c0",-- 12
x"00000",-- 0
x"fff40",-- -12
x"fffe0",-- -2
x"00390",-- 57
x"005d0",-- 93
x"001c0",-- 28
x"ffd50",-- -43
x"ffea0",-- -22
x"001b0",-- 27
x"00210",-- 33
x"00120",-- 18
x"00250",-- 37
x"002f0",-- 47
x"00250",-- 37
x"00020",-- 2
x"ffe50",-- -27
x"fffd0",-- -3
x"000a0",-- 10
x"ffee0",-- -18
x"ffc60",-- -58
x"ffd50",-- -43
x"fff90",-- -7
x"ffee0",-- -18
x"ffc60",-- -58
x"ffb80",-- -72
x"ff950",-- -107
x"ff8f0",-- -113
x"ffad0",-- -83
x"ffad0",-- -83
x"ffb80",-- -72
x"ffcc0",-- -52
x"ffd80",-- -40
x"ffe00",-- -32
x"00000",-- 0
x"00000",-- 0
x"ffe20",-- -30
x"ffce0",-- -50
x"fffb0",-- -5
x"001e0",-- 30
x"00160",-- 22
x"00030",-- 3
x"00000",-- 0
x"00000",-- 0
x"fffd0",-- -3
x"00000",-- 0
x"00070",-- 7
x"00020",-- 2
x"00000",-- 0
x"00050",-- 5
x"fff60",-- -10
x"ffec0",-- -20
x"fff10",-- -15
x"ffe90",-- -23
x"ffd80",-- -40
x"ffea0",-- -22
x"fff40",-- -12
x"000f0",-- 15
x"00110",-- 17
x"00160",-- 22
x"00250",-- 37
x"00080",-- 8
x"00080",-- 8
x"00370",-- 55
x"00640",-- 100
x"004b0",-- 75
x"00370",-- 55
x"003e0",-- 62
x"005f0",-- 95
x"007d0",-- 125
x"006c0",-- 108
x"00410",-- 65
x"00250",-- 37
x"002a0",-- 42
x"00250",-- 37
x"00120",-- 18
x"00080",-- 8
x"00020",-- 2
x"000c0",-- 12
x"fffb0",-- -5
x"00020",-- 2
x"00280",-- 40
x"00250",-- 37
x"fff60",-- -10
x"ffc20",-- -62
x"ffe50",-- -27
x"00140",-- 20
x"002f0",-- 47
x"00230",-- 35
x"fff40",-- -12
x"ffe50",-- -27
x"ffdd0",-- -35
x"ffee0",-- -18
x"fffe0",-- -2
x"fffb0",-- -5
x"00020",-- 2
x"fff80",-- -8
x"fff30",-- -13
x"00000",-- 0
x"00020",-- 2
x"ffe90",-- -23
x"ffc60",-- -58
x"ffd50",-- -43
x"ffe40",-- -28
x"fff40",-- -12
x"fffb0",-- -5
x"000c0",-- 12
x"00160",-- 22
x"00000",-- 0
x"000f0",-- 15
x"001b0",-- 27
x"00170",-- 23
x"000c0",-- 12
x"ffe90",-- -23
x"ffce0",-- -50
x"ffee0",-- -18
x"00160",-- 22
x"00320",-- 50
x"00280",-- 40
x"fff40",-- -12
x"ffce0",-- -50
x"ffee0",-- -18
x"002b0",-- 43
x"00410",-- 65
x"002b0",-- 43
x"fffe0",-- -2
x"00000",-- 0
x"00070",-- 7
x"00020",-- 2
x"fff80",-- -8
x"fff10",-- -15
x"00080",-- 8
x"000f0",-- 15
x"000f0",-- 15
x"fff40",-- -12
x"ffea0",-- -22
x"fff40",-- -12
x"000a0",-- 10
x"00250",-- 37
x"00190",-- 25
x"fff60",-- -10
x"ffe20",-- -30
x"000f0",-- 15
x"00370",-- 55
x"00000",-- 0
x"ffb50",-- -75
x"ffb50",-- -75
x"ffec0",-- -20
x"00190",-- 25
x"00120",-- 18
x"ffd80",-- -40
x"ffab0",-- -85
x"ffc90",-- -55
x"00080",-- 8
x"004b0",-- 75
x"00520",-- 82
x"002b0",-- 43
x"fff40",-- -12
x"fff10",-- -15
x"00250",-- 37
x"00500",-- 80
x"002a0",-- 42
x"fffb0",-- -5
x"ffe90",-- -23
x"00000",-- 0
x"00120",-- 18
x"fffd0",-- -3
x"ffea0",-- -22
x"ffd80",-- -40
x"ffe20",-- -30
x"fff60",-- -10
x"fff80",-- -8
x"ffe20",-- -30
x"ffc90",-- -55
x"ffdd0",-- -35
x"fff40",-- -12
x"fffe0",-- -2
x"fff90",-- -7
x"ffc60",-- -58
x"ffb50",-- -75
x"ffe20",-- -30
x"002b0",-- 43
x"00320",-- 50
x"000c0",-- 12
x"fff90",-- -7
x"fffe0",-- -2
x"00140",-- 20
x"00260",-- 38
x"001c0",-- 28
x"fffd0",-- -3
x"00080",-- 8
x"001b0",-- 27
x"00000",-- 0
x"ffc20",-- -62
x"ffc90",-- -55
x"00020",-- 2
x"00020",-- 2
x"ffd80",-- -40
x"ffc10",-- -63
x"ffc90",-- -55
x"fffd0",-- -3
x"00210",-- 33
x"ffef0",-- -17
x"ff950",-- -107
x"ff860",-- -122
x"ffd50",-- -43
x"00170",-- 23
x"fffe0",-- -2
x"ffbf0",-- -65
x"ffb20",-- -78
x"ffd00",-- -48
x"00000",-- 0
x"001b0",-- 27
x"00110",-- 17
x"00050",-- 5
x"00000",-- 0
x"00000",-- 0
x"00080",-- 8
x"000a0",-- 10
x"00000",-- 0
x"ffb00",-- -80
x"ff7c0",-- -132
x"ff9e0",-- -98
x"ffdb0",-- -37
x"00080",-- 8
x"00000",-- 0
x"ffd30",-- -45
x"ffb70",-- -73
x"ffb80",-- -72
x"ffb70",-- -73
x"ffb20",-- -78
x"ffd50",-- -43
x"ffd10",-- -47
x"ffbd0",-- -67
x"ffc10",-- -63
x"ffe50",-- -27
x"ffdf0",-- -33
x"ffdd0",-- -35
x"ffea0",-- -22
x"ffdf0",-- -33
x"00000",-- 0
x"00230",-- 35
x"000f0",-- 15
x"ffee0",-- -18
x"ffda0",-- -38
x"ffe20",-- -30
x"ffe20",-- -30
x"ffc70",-- -57
x"ffc10",-- -63
x"ffa90",-- -87
x"ff9f0",-- -97
x"ffa10",-- -95
x"ffc40",-- -60
x"ffe50",-- -27
x"ffd80",-- -40
x"ffa30",-- -93
x"ff860",-- -122
x"ffb00",-- -80
x"ffe20",-- -30
x"ffe50",-- -27
x"ff9c0",-- -100
x"ff680",-- -152
x"ff950",-- -107
x"fff40",-- -12
x"00170",-- 23
x"ffe20",-- -30
x"ff970",-- -105
x"ff900",-- -112
x"ffbf0",-- -65
x"fffd0",-- -3
x"000f0",-- 15
x"ffee0",-- -18
x"ffbf0",-- -65
x"ffb20",-- -78
x"ffb20",-- -78
x"ffd10",-- -47
x"fff10",-- -15
x"ffd30",-- -45
x"ff990",-- -103
x"ff9f0",-- -97
x"ffd60",-- -42
x"ffe20",-- -30
x"ffcb0",-- -53
x"ffc90",-- -55
x"ffce0",-- -50
x"ffd00",-- -48
x"ffd00",-- -48
x"ffc90",-- -55
x"ffdb0",-- -37
x"ffe20",-- -30
x"ffdb0",-- -37
x"ffc10",-- -63
x"ffdb0",-- -37
x"fff80",-- -8
x"ffd50",-- -43
x"ffc60",-- -58
x"ffdf0",-- -33
x"fffb0",-- -5
x"ffe70",-- -25
x"ffc20",-- -62
x"ff860",-- -122
x"ff970",-- -105
x"ffe20",-- -30
x"ffea0",-- -22
x"ff990",-- -103
x"ff900",-- -112
x"fffe0",-- -2
x"00410",-- 65
x"00160",-- 22
x"ffc90",-- -55
x"ff9c0",-- -100
x"ffb30",-- -77
x"00110",-- 17
x"00410",-- 65
x"00160",-- 22
x"ffda0",-- -38
x"ffd80",-- -40
x"001b0",-- 27
x"005a0",-- 90
x"00350",-- 53
x"ffd10",-- -47
x"ffb30",-- -77
x"ffea0",-- -22
x"000f0",-- 15
x"00000",-- 0
x"fffb0",-- -5
x"00000",-- 0
x"00020",-- 2
x"ffe50",-- -27
x"ffdb0",-- -37
x"fff10",-- -15
x"00020",-- 2
x"fff90",-- -7
x"ffdd0",-- -35
x"ffd10",-- -47
x"ffdb0",-- -37
x"fff30",-- -13
x"fffe0",-- -2
x"fff60",-- -10
x"ffc90",-- -55
x"ffa80",-- -88
x"ffbc0",-- -68
x"ffea0",-- -22
x"fffd0",-- -3
x"ffea0",-- -22
x"ffc90",-- -55
x"ffbf0",-- -65
x"ffd60",-- -42
x"00000",-- 0
x"00000",-- 0
x"fff40",-- -12
x"ffe70",-- -25
x"fff10",-- -15
x"fffb0",-- -5
x"00030",-- 3
x"00320",-- 50
x"002a0",-- 42
x"000d0",-- 13
x"00050",-- 5
x"000c0",-- 12
x"00020",-- 2
x"ffee0",-- -18
x"ffec0",-- -20
x"ffee0",-- -18
x"fff90",-- -7
x"fff40",-- -12
x"ffdf0",-- -33
x"ffdd0",-- -35
x"00070",-- 7
x"003e0",-- 62
x"002f0",-- 47
x"00020",-- 2
x"ffee0",-- -18
x"ffdd0",-- -35
x"ffee0",-- -18
x"00160",-- 22
x"001b0",-- 27
x"000d0",-- 13
x"001c0",-- 28
x"00210",-- 33
x"00030",-- 3
x"000f0",-- 15
x"002b0",-- 43
x"000c0",-- 12
x"00000",-- 0
x"000c0",-- 12
x"000f0",-- 15
x"00110",-- 17
x"00250",-- 37
x"000d0",-- 13
x"ffe90",-- -23
x"ffdf0",-- -33
x"ffd10",-- -47
x"ffb50",-- -75
x"ffb70",-- -73
x"ffdb0",-- -37
x"ffe50",-- -27
x"ffee0",-- -18
x"ffe50",-- -27
x"ffe50",-- -27
x"ffea0",-- -22
x"fffe0",-- -2
x"00000",-- 0
x"ffe90",-- -23
x"ffe50",-- -27
x"fff10",-- -15
x"00000",-- 0
x"00000",-- 0
x"00120",-- 18
x"001b0",-- 27
x"00120",-- 18
x"00120",-- 18
x"00250",-- 37
x"00320",-- 50
x"00260",-- 38
x"00350",-- 53
x"002d0",-- 45
x"00160",-- 22
x"00020",-- 2
x"00030",-- 3
x"00050",-- 5
x"00030",-- 3
x"00320",-- 50
x"003a0",-- 58
x"001c0",-- 28
x"00030",-- 3
x"00050",-- 5
x"00140",-- 20
x"003a0",-- 58
x"00480",-- 72
x"002b0",-- 43
x"00230",-- 35
x"00190",-- 25
x"00250",-- 37
x"002f0",-- 47
x"002f0",-- 47
x"00320",-- 50
x"00280",-- 40
x"00320",-- 50
x"00230",-- 35
x"00190",-- 25
x"002f0",-- 47
x"003e0",-- 62
x"003e0",-- 62
x"00190",-- 25
x"fff90",-- -7
x"ffef0",-- -17
x"00050",-- 5
x"00300",-- 48
x"00370",-- 55
x"00000",-- 0
x"ffee0",-- -18
x"fff80",-- -8
x"00000",-- 0
x"000f0",-- 15
x"002b0",-- 43
x"001b0",-- 27
x"00050",-- 5
x"001b0",-- 27
x"00430",-- 67
x"00570",-- 87
x"00570",-- 87
x"003e0",-- 62
x"001b0",-- 27
x"000d0",-- 13
x"000f0",-- 15
x"00070",-- 7
x"00020",-- 2
x"00120",-- 18
x"00210",-- 33
x"000c0",-- 12
x"fff10",-- -15
x"fffd0",-- -3
x"000f0",-- 15
x"000c0",-- 12
x"fffd0",-- -3
x"00050",-- 5
x"00080",-- 8
x"00020",-- 2
x"000c0",-- 12
x"00370",-- 55
x"00610",-- 97
x"005f0",-- 95
x"002f0",-- 47
x"00050",-- 5
x"00160",-- 22
x"004e0",-- 78
x"00780",-- 120
x"00410",-- 65
x"ffe20",-- -30
x"ffbc0",-- -68
x"fff10",-- -15
x"002d0",-- 45
x"00250",-- 37
x"ffd10",-- -47
x"ff920",-- -110
x"ff850",-- -123
x"ffc90",-- -55
x"fffb0",-- -5
x"ffd50",-- -43
x"ffa90",-- -87
x"ff8a0",-- -118
x"ffa90",-- -87
x"ffd80",-- -40
x"fffe0",-- -2
x"fff40",-- -12
x"ffda0",-- -38
x"ffc90",-- -55
x"ffdf0",-- -33
x"000f0",-- 15
x"00370",-- 55
x"00280",-- 40
x"00250",-- 37
x"00300",-- 48
x"001b0",-- 27
x"00160",-- 22
x"00050",-- 5
x"00070",-- 7
x"00080",-- 8
x"000d0",-- 13
x"000f0",-- 15
x"000a0",-- 10
x"00030",-- 3
x"ffe70",-- -25
x"ffe50",-- -27
x"ffe50",-- -27
x"ffdb0",-- -37
x"ffd10",-- -47
x"ffdb0",-- -37
x"ffee0",-- -18
x"fff80",-- -8
x"fff30",-- -13
x"ffe20",-- -30
x"fff80",-- -8
x"001b0",-- 27
x"00200",-- 32
x"00000",-- 0
x"fff10",-- -15
x"00070",-- 7
x"00280",-- 40
x"003e0",-- 62
x"00410",-- 65
x"00230",-- 35
x"00000",-- 0
x"00050",-- 5
x"002a0",-- 42
x"002b0",-- 43
x"fff10",-- -15
x"ffb50",-- -75
x"ffbf0",-- -65
x"ffea0",-- -22
x"00000",-- 0
x"ffe90",-- -23
x"ffab0",-- -85
x"ffb70",-- -73
x"ffe90",-- -23
x"fff80",-- -8
x"ffe50",-- -27
x"ffda0",-- -38
x"ffe00",-- -32
x"00030",-- 3
x"00440",-- 68
x"00410",-- 65
x"000c0",-- 12
x"fff80",-- -8
x"000c0",-- 12
x"002d0",-- 45
x"003c0",-- 60
x"00410",-- 65
x"00160",-- 22
x"00000",-- 0
x"001b0",-- 27
x"002f0",-- 47
x"00320",-- 50
x"00260",-- 38
x"00120",-- 18
x"ffea0",-- -22
x"ffdb0",-- -37
x"fffe0",-- -2
x"00020",-- 2
x"fffe0",-- -2
x"fffb0",-- -5
x"fffb0",-- -5
x"ffe70",-- -25
x"ffdb0",-- -37
x"ffec0",-- -20
x"00030",-- 3
x"00080",-- 8
x"00050",-- 5
x"00000",-- 0
x"ffe90",-- -23
x"ffe50",-- -27
x"fffb0",-- -5
x"00070",-- 7
x"00120",-- 18
x"000f0",-- 15
x"fffe0",-- -2
x"fffb0",-- -5
x"00000",-- 0
x"001b0",-- 27
x"00000",-- 0
x"ffe90",-- -23
x"ffd50",-- -43
x"ffc20",-- -62
x"ffdb0",-- -37
x"ffe40",-- -28
x"ffdf0",-- -33
x"ffdf0",-- -33
x"00020",-- 2
x"00070",-- 7
x"ffee0",-- -18
x"ffe40",-- -28
x"00080",-- 8
x"002f0",-- 47
x"00370",-- 55
x"00370",-- 55
x"000c0",-- 12
x"00000",-- 0
x"00160",-- 22
x"001e0",-- 30
x"000c0",-- 12
x"00050",-- 5
x"00020",-- 2
x"000c0",-- 12
x"002f0",-- 47
x"002b0",-- 43
x"fff10",-- -15
x"ffc90",-- -55
x"ffe00",-- -32
x"fffb0",-- -5
x"fff40",-- -12
x"ffd00",-- -48
x"ffd50",-- -43
x"fff40",-- -12
x"000f0",-- 15
x"00080",-- 8
x"ffdd0",-- -35
x"ffe70",-- -25
x"000f0",-- 15
x"001c0",-- 28
x"000a0",-- 10
x"ffea0",-- -22
x"ffdb0",-- -37
x"ffe00",-- -32
x"fffd0",-- -3
x"fffd0",-- -3
x"ffd10",-- -47
x"ffba0",-- -70
x"ffc20",-- -62
x"ffd60",-- -42
x"ffe40",-- -28
x"fff60",-- -10
x"00000",-- 0
x"ffe90",-- -23
x"ffdb0",-- -37
x"ffdb0",-- -37
x"ffc90",-- -55
x"ffef0",-- -17
x"00140",-- 20
x"00170",-- 23
x"ffec0",-- -20
x"ffc60",-- -58
x"ffd30",-- -45
x"fffe0",-- -2
x"00250",-- 37
x"fff80",-- -8
x"ffbd0",-- -67
x"ffce0",-- -50
x"fff80",-- -8
x"000d0",-- 13
x"000a0",-- 10
x"ffec0",-- -20
x"ffec0",-- -20
x"000f0",-- 15
x"001b0",-- 27
x"00080",-- 8
x"fff40",-- -12
x"ffe40",-- -28
x"fffb0",-- -5
x"000f0",-- 15
x"00170",-- 23
x"fff40",-- -12
x"ffda0",-- -38
x"fffd0",-- -3
x"00170",-- 23
x"00140",-- 20
x"00000",-- 0
x"ffef0",-- -17
x"fff60",-- -10
x"00000",-- 0
x"fffb0",-- -5
x"ffdd0",-- -35
x"ffd50",-- -43
x"ffdb0",-- -37
x"ffc20",-- -62
x"ffc10",-- -63
x"ffc60",-- -58
x"ffdb0",-- -37
x"ffee0",-- -18
x"ffe00",-- -32
x"ffc20",-- -62
x"ffc20",-- -62
x"ffe70",-- -25
x"ffec0",-- -20
x"ffbd0",-- -67
x"ff9c0",-- -100
x"ff990",-- -103
x"ffa10",-- -95
x"ffb30",-- -77
x"ffba0",-- -70
x"ffc90",-- -55
x"ffd50",-- -43
x"ffc60",-- -58
x"ffc60",-- -58
x"ffe00",-- -32
x"ffe90",-- -23
x"ffd60",-- -42
x"ffce0",-- -50
x"ffbd0",-- -67
x"ffc10",-- -63
x"ffc60",-- -58
x"ffc90",-- -55
x"ffb50",-- -75
x"ffa90",-- -87
x"ff9a0",-- -102
x"ff8a0",-- -118
x"ffa10",-- -95
x"ffce0",-- -50
x"ffe40",-- -28
x"ffd00",-- -48
x"ffbd0",-- -67
x"ffbd0",-- -67
x"ffe50",-- -27
x"fffb0",-- -5
x"fff80",-- -8
x"ffc40",-- -60
x"ffae0",-- -82
x"ffce0",-- -50
x"fff30",-- -13
x"000f0",-- 15
x"00170",-- 23
x"00110",-- 17
x"fff80",-- -8
x"fff80",-- -8
x"ffe20",-- -30
x"ffdd0",-- -35
x"fff80",-- -8
x"00000",-- 0
x"00000",-- 0
x"fff60",-- -10
x"ffea0",-- -22
x"ffee0",-- -18
x"fffe0",-- -2
x"fff80",-- -8
x"ffdf0",-- -33
x"ffd50",-- -43
x"ffd10",-- -47
x"ffd80",-- -40
x"ffe70",-- -25
x"00000",-- 0
x"fff80",-- -8
x"ffc60",-- -58
x"ffab0",-- -85
x"ffb50",-- -75
x"ffd30",-- -45
x"ffcc0",-- -52
x"ffad0",-- -83
x"ff850",-- -123
x"ff810",-- -127
x"ff970",-- -105
x"ffb50",-- -75
x"ffb70",-- -73
x"ffc70",-- -57
x"ffdb0",-- -37
x"ffc40",-- -60
x"ffad0",-- -83
x"ffb70",-- -73
x"fff40",-- -12
x"00120",-- 18
x"00080",-- 8
x"ffec0",-- -20
x"ffd10",-- -47
x"ffe50",-- -27
x"000a0",-- 10
x"001b0",-- 27
x"00250",-- 37
x"00080",-- 8
x"ffe70",-- -25
x"ffee0",-- -18
x"000f0",-- 15
x"002b0",-- 43
x"00280",-- 40
x"00050",-- 5
x"00000",-- 0
x"00000",-- 0
x"00030",-- 3
x"fffb0",-- -5
x"fff40",-- -12
x"00050",-- 5
x"00000",-- 0
x"fff10",-- -15
x"ffee0",-- -18
x"fffd0",-- -3
x"000a0",-- 10
x"00120",-- 18
x"000f0",-- 15
x"00080",-- 8
x"000c0",-- 12
x"00000",-- 0
x"ffe50",-- -27
x"fff10",-- -15
x"00080",-- 8
x"00160",-- 22
x"000f0",-- 15
x"fff80",-- -8
x"ffdd0",-- -35
x"fff10",-- -15
x"00160",-- 22
x"00160",-- 22
x"00050",-- 5
x"00070",-- 7
x"00120",-- 18
x"00230",-- 35
x"00230",-- 35
x"001e0",-- 30
x"00120",-- 18
x"00250",-- 37
x"00280",-- 40
x"00170",-- 23
x"00080",-- 8
x"00000",-- 0
x"00020",-- 2
x"fffe0",-- -2
x"ffec0",-- -20
x"ffdd0",-- -35
x"ffd80",-- -40
x"ffe90",-- -23
x"fff10",-- -15
x"ffe00",-- -32
x"ffd30",-- -45
x"ffc60",-- -58
x"ffc60",-- -58
x"ffbf0",-- -65
x"ffc60",-- -58
x"ffdb0",-- -37
x"ffd80",-- -40
x"ffc10",-- -63
x"ffc60",-- -58
x"ffdf0",-- -33
x"ffea0",-- -22
x"fff80",-- -8
x"fffd0",-- -3
x"ffe40",-- -28
x"ffcb0",-- -53
x"ffd10",-- -47
x"ffd60",-- -42
x"fff10",-- -15
x"fffe0",-- -2
x"ffea0",-- -22
x"ffe50",-- -27
x"ffe50",-- -27
x"ffef0",-- -17
x"ffdb0",-- -37
x"ffc60",-- -58
x"ffd80",-- -40
x"fff80",-- -8
x"fff60",-- -10
x"ffdf0",-- -33
x"ffc20",-- -62
x"ffc90",-- -55
x"fffb0",-- -5
x"00000",-- 0
x"ffdf0",-- -33
x"ffcc0",-- -52
x"ffe50",-- -27
x"00140",-- 20
x"002d0",-- 45
x"002a0",-- 42
x"001b0",-- 27
x"000f0",-- 15
x"00140",-- 20
x"000c0",-- 12
x"00120",-- 18
x"00000",-- 0
x"ffee0",-- -18
x"ffee0",-- -18
x"fffb0",-- -5
x"001b0",-- 27
x"002a0",-- 42
x"00140",-- 20
x"fff80",-- -8
x"fffe0",-- -2
x"00020",-- 2
x"00080",-- 8
x"000f0",-- 15
x"00080",-- 8
x"00000",-- 0
x"fff40",-- -12
x"fff80",-- -8
x"00000",-- 0
x"000a0",-- 10
x"000c0",-- 12
x"00020",-- 2
x"00000",-- 0
x"00110",-- 17
x"00200",-- 32
x"00280",-- 40
x"00260",-- 38
x"00320",-- 50
x"002b0",-- 43
x"002b0",-- 43
x"00110",-- 17
x"fffd0",-- -3
x"00030",-- 3
x"00000",-- 0
x"ffee0",-- -18
x"ffdf0",-- -33
x"ffdd0",-- -35
x"ffdb0",-- -37
x"fffb0",-- -5
x"001b0",-- 27
x"001e0",-- 30
x"000a0",-- 10
x"fff10",-- -15
x"ffea0",-- -22
x"fff80",-- -8
x"00120",-- 18
x"00160",-- 22
x"00000",-- 0
x"ffea0",-- -22
x"ffe40",-- -28
x"00120",-- 18
x"003c0",-- 60
x"00460",-- 70
x"002d0",-- 45
x"00110",-- 17
x"00080",-- 8
x"00140",-- 20
x"00370",-- 55
x"003c0",-- 60
x"001e0",-- 30
x"000c0",-- 12
x"ffdf0",-- -33
x"ffc40",-- -60
x"ffcc0",-- -52
x"ffdd0",-- -35
x"fffd0",-- -3
x"fff60",-- -10
x"ffd60",-- -42
x"ffb70",-- -73
x"ffd50",-- -43
x"00160",-- 22
x"001e0",-- 30
x"fff40",-- -12
x"ffd10",-- -47
x"ffe20",-- -30
x"00000",-- 0
x"00030",-- 3
x"00030",-- 3
x"00000",-- 0
x"00020",-- 2
x"000f0",-- 15
x"00210",-- 33
x"003f0",-- 63
x"00440",-- 68
x"00280",-- 40
x"001e0",-- 30
x"001b0",-- 27
x"00250",-- 37
x"00390",-- 57
x"001c0",-- 28
x"fffb0",-- -5
x"fff60",-- -10
x"fff90",-- -7
x"00000",-- 0
x"00190",-- 25
x"001e0",-- 30
x"00000",-- 0
x"ffd00",-- -48
x"ffb80",-- -72
x"ffec0",-- -20
x"000a0",-- 10
x"00020",-- 2
x"ffce0",-- -50
x"ffb30",-- -77
x"ffdf0",-- -33
x"002f0",-- 47
x"00530",-- 83
x"00230",-- 35
x"fff90",-- -7
x"ffdf0",-- -33
x"00080",-- 8
x"003a0",-- 58
x"002f0",-- 47
x"00000",-- 0
x"ffe00",-- -32
x"ffe20",-- -30
x"00000",-- 0
x"00200",-- 32
x"00070",-- 7
x"ffdb0",-- -37
x"ffd80",-- -40
x"ffe20",-- -30
x"00000",-- 0
x"00190",-- 25
x"00050",-- 5
x"fff10",-- -15
x"ffe90",-- -23
x"fff30",-- -13
x"fff60",-- -10
x"fff10",-- -15
x"fff90",-- -7
x"fff80",-- -8
x"fff10",-- -15
x"ffea0",-- -22
x"ffe90",-- -23
x"ffe20",-- -30
x"fff30",-- -13
x"00000",-- 0
x"00000",-- 0
x"fffe0",-- -2
x"fff60",-- -10
x"00000",-- 0
x"00000",-- 0
x"fffd0",-- -3
x"00080",-- 8
x"00190",-- 25
x"00280",-- 40
x"00320",-- 50
x"00080",-- 8
x"ffee0",-- -18
x"fff90",-- -7
x"00140",-- 20
x"000d0",-- 13
x"ffee0",-- -18
x"ffda0",-- -38
x"ffe20",-- -30
x"000c0",-- 12
x"00250",-- 37
x"00020",-- 2
x"ffd50",-- -43
x"ffd00",-- -48
x"ffef0",-- -17
x"00050",-- 5
x"ffdf0",-- -33
x"ffb00",-- -80
x"ffbf0",-- -65
x"fffd0",-- -3
x"002f0",-- 47
x"001e0",-- 30
x"fffd0",-- -3
x"00000",-- 0
x"00280",-- 40
x"00340",-- 52
x"00120",-- 18
x"ffdb0",-- -37
x"ffe20",-- -30
x"00030",-- 3
x"002f0",-- 47
x"002a0",-- 42
x"fff80",-- -8
x"ffce0",-- -50
x"ffcb0",-- -53
x"ffe00",-- -32
x"fff10",-- -15
x"ffee0",-- -18
x"ffd80",-- -40
x"ffcc0",-- -52
x"ffd60",-- -42
x"00020",-- 2
x"000f0",-- 15
x"fffd0",-- -3
x"fff40",-- -12
x"00000",-- 0
x"00210",-- 33
x"004b0",-- 75
x"00500",-- 80
x"00340",-- 52
x"00350",-- 53
x"004e0",-- 78
x"005c0",-- 92
x"00440",-- 68
x"00260",-- 38
x"00160",-- 22
x"00250",-- 37
x"002f0",-- 47
x"001e0",-- 30
x"00050",-- 5
x"fff40",-- -12
x"00000",-- 0
x"000f0",-- 15
x"000a0",-- 10
x"fff10",-- -15
x"fff80",-- -8
x"000c0",-- 12
x"000f0",-- 15
x"fff60",-- -10
x"ffec0",-- -20
x"ffea0",-- -22
x"00030",-- 3
x"00250",-- 37
x"00120",-- 18
x"00050",-- 5
x"000f0",-- 15
x"002f0",-- 47
x"002f0",-- 47
x"000f0",-- 15
x"fffe0",-- -2
x"00000",-- 0
x"00260",-- 38
x"00480",-- 72
x"00210",-- 33
x"ffee0",-- -18
x"ffe50",-- -27
x"00160",-- 22
x"00440",-- 68
x"00250",-- 37
x"ffe90",-- -23
x"ffda0",-- -38
x"00120",-- 18
x"004e0",-- 78
x"004b0",-- 75
x"00020",-- 2
x"ffd10",-- -47
x"ffe90",-- -23
x"001b0",-- 27
x"00350",-- 53
x"00000",-- 0
x"ffce0",-- -50
x"ffc20",-- -62
x"fff80",-- -8
x"00160",-- 22
x"fff90",-- -7
x"ffd10",-- -47
x"ffb80",-- -72
x"ffcb0",-- -53
x"ffef0",-- -17
x"fffe0",-- -2
x"ffec0",-- -20
x"ffdd0",-- -35
x"ffea0",-- -22
x"fffb0",-- -5
x"fffb0",-- -5
x"ffec0",-- -20
x"ffea0",-- -22
x"00000",-- 0
x"00160",-- 22
x"00050",-- 5
x"fff80",-- -8
x"00000",-- 0
x"00160",-- 22
x"00000",-- 0
x"ffe00",-- -32
x"ffb50",-- -75
x"ffb80",-- -72
x"ffe50",-- -27
x"fff80",-- -8
x"fff60",-- -10
x"ffd30",-- -45
x"ffba0",-- -70
x"ffb00",-- -80
x"ffbf0",-- -65
x"ffb80",-- -72
x"ffb20",-- -78
x"ffbc0",-- -68
x"ffd10",-- -47
x"ffdd0",-- -35
x"ffdb0",-- -37
x"ffd50",-- -43
x"ffe90",-- -23
x"fff40",-- -12
x"ffec0",-- -20
x"ffdb0",-- -37
x"ffda0",-- -38
x"fffe0",-- -2
x"000d0",-- 13
x"00050",-- 5
x"ffea0",-- -22
x"ffdf0",-- -33
x"fff60",-- -10
x"001e0",-- 30
x"00190",-- 25
x"fffd0",-- -3
x"ffdb0",-- -37
x"ffd80",-- -40
x"fff80",-- -8
x"00020",-- 2
x"fffb0",-- -5
x"ffc60",-- -58
x"ffa60",-- -90
x"ffbf0",-- -65
x"00000",-- 0
x"001e0",-- 30
x"00120",-- 18
x"ffee0",-- -18
x"ffb50",-- -75
x"ffb70",-- -73
x"ffdf0",-- -33
x"000d0",-- 13
x"001b0",-- 27
x"fff80",-- -8
x"ffe50",-- -27
x"ffdf0",-- -33
x"ffdf0",-- -33
x"fff30",-- -13
x"fff10",-- -15
x"ffe40",-- -28
x"ffc60",-- -58
x"ffb20",-- -78
x"ffd00",-- -48
x"ffea0",-- -22
x"00080",-- 8
x"fff90",-- -7
x"ffb20",-- -78
x"ffa30",-- -93
x"ffbc0",-- -68
x"fff10",-- -15
x"00000",-- 0
x"ffd80",-- -40
x"ff950",-- -107
x"ff8d0",-- -115
x"ffdd0",-- -35
x"00210",-- 33
x"00140",-- 20
x"ffd80",-- -40
x"ff9e0",-- -98
x"ffb20",-- -78
x"fffe0",-- -2
x"001e0",-- 30
x"fffb0",-- -5
x"ffb80",-- -72
x"ff9f0",-- -97
x"ffc90",-- -55
x"00050",-- 5
x"00230",-- 35
x"00000",-- 0
x"ffdb0",-- -37
x"ffe20",-- -30
x"ffea0",-- -22
x"fff30",-- -13
x"fff60",-- -10
x"fff10",-- -15
x"fff10",-- -15
x"ffef0",-- -17
x"ffd60",-- -42
x"ffc60",-- -58
x"ffd30",-- -45
x"ffef0",-- -17
x"00000",-- 0
x"fff40",-- -12
x"ffe20",-- -30
x"ffd60",-- -42
x"ffdf0",-- -33
x"fffb0",-- -5
x"00000",-- 0
x"00140",-- 20
x"00080",-- 8
x"ffd80",-- -40
x"ffc70",-- -57
x"ffea0",-- -22
x"001b0",-- 27
x"00320",-- 50
x"00030",-- 3
x"ffce0",-- -50
x"ffd30",-- -45
x"00000",-- 0
x"00250",-- 37
x"00190",-- 25
x"ffe40",-- -28
x"ffbc0",-- -68
x"ffc10",-- -63
x"ffdf0",-- -33
x"fff80",-- -8
x"fff10",-- -15
x"ffd00",-- -48
x"ffb30",-- -77
x"ffbf0",-- -65
x"ffe40",-- -28
x"00110",-- 17
x"00280",-- 40
x"00120",-- 18
x"ffee0",-- -18
x"ffe20",-- -30
x"fff10",-- -15
x"001e0",-- 30
x"00370",-- 55
x"001e0",-- 30
x"fff90",-- -7
x"ffc10",-- -63
x"ffd10",-- -47
x"00070",-- 7
x"00120",-- 18
x"fff10",-- -15
x"ffbc0",-- -68
x"ffa90",-- -87
x"ffd50",-- -43
x"fff90",-- -7
x"ffea0",-- -22
x"ffc70",-- -57
x"ffa30",-- -93
x"ffc90",-- -55
x"00000",-- 0
x"fffe0",-- -2
x"ffdd0",-- -35
x"ffc70",-- -57
x"ffd30",-- -45
x"00000",-- 0
x"00080",-- 8
x"ffe50",-- -27
x"ffc20",-- -62
x"ffa90",-- -87
x"ffc90",-- -55
x"fff40",-- -12
x"00050",-- 5
x"fffd0",-- -3
x"ffe90",-- -23
x"ffd10",-- -47
x"ffdf0",-- -33
x"fff80",-- -8
x"ffea0",-- -22
x"ffe70",-- -25
x"ffdd0",-- -35
x"ffdf0",-- -33
x"ffe90",-- -23
x"fff30",-- -13
x"ffef0",-- -17
x"fff40",-- -12
x"fffb0",-- -5
x"ffdb0",-- -37
x"ffc70",-- -57
x"ffd30",-- -45
x"00000",-- 0
x"000f0",-- 15
x"fff90",-- -7
x"ffc90",-- -55
x"ffa40",-- -92
x"ffb20",-- -78
x"ffce0",-- -50
x"ffe20",-- -30
x"ffc70",-- -57
x"ffa30",-- -93
x"ff9a0",-- -102
x"ffb30",-- -77
x"ffdb0",-- -37
x"ffef0",-- -17
x"ffea0",-- -22
x"ffd10",-- -47
x"ffce0",-- -50
x"ffdf0",-- -33
x"fff30",-- -13
x"fffb0",-- -5
x"00000",-- 0
x"fff10",-- -15
x"ffee0",-- -18
x"fff10",-- -15
x"fff40",-- -12
x"00000",-- 0
x"00110",-- 17
x"00190",-- 25
x"00000",-- 0
x"fffb0",-- -5
x"00020",-- 2
x"001c0",-- 28
x"00390",-- 57
x"001e0",-- 30
x"fff40",-- -12
x"ffd50",-- -43
x"ffdb0",-- -37
x"fffb0",-- -5
x"00140",-- 20
x"00070",-- 7
x"ffe90",-- -23
x"ffce0",-- -50
x"ffdb0",-- -37
x"00030",-- 3
x"001e0",-- 30
x"000a0",-- 10
x"fff10",-- -15
x"ffe50",-- -27
x"ffe70",-- -25
x"000c0",-- 12
x"00110",-- 17
x"00080",-- 8
x"fffb0",-- -5
x"fffb0",-- -5
x"00000",-- 0
x"fffb0",-- -5
x"fff80",-- -8
x"fffb0",-- -5
x"00000",-- 0
x"fff90",-- -7
x"ffe20",-- -30
x"ffd80",-- -40
x"ffec0",-- -20
x"fff80",-- -8
x"fffe0",-- -2
x"fff40",-- -12
x"ffdb0",-- -37
x"ffd50",-- -43
x"ffe40",-- -28
x"fff80",-- -8
x"00000",-- 0
x"fffb0",-- -5
x"ffe70",-- -25
x"fff10",-- -15
x"ffee0",-- -18
x"00000",-- 0
x"00030",-- 3
x"00000",-- 0
x"fffb0",-- -5
x"ffef0",-- -17
x"fff10",-- -15
x"ffef0",-- -17
x"fff10",-- -15
x"ffe90",-- -23
x"fff10",-- -15
x"fff60",-- -10
x"ffea0",-- -22
x"ffe50",-- -27
x"fff10",-- -15
x"00000",-- 0
x"fff80",-- -8
x"ffea0",-- -22
x"ffe70",-- -25
x"fff80",-- -8
x"fffb0",-- -5
x"00000",-- 0
x"00020",-- 2
x"fffb0",-- -5
x"00000",-- 0
x"000f0",-- 15
x"001b0",-- 27
x"00230",-- 35
x"001e0",-- 30
x"000c0",-- 12
x"00000",-- 0
x"00000",-- 0
x"000f0",-- 15
x"00120",-- 18
x"000a0",-- 10
x"fff40",-- -12
x"ffe90",-- -23
x"00000",-- 0
x"000f0",-- 15
x"001b0",-- 27
x"00190",-- 25
x"fff60",-- -10
x"ffec0",-- -20
x"fff30",-- -13
x"00000",-- 0
x"fffe0",-- -2
x"fff40",-- -12
x"ffe40",-- -28
x"ffdb0",-- -37
x"ffea0",-- -22
x"fff10",-- -15
x"fff30",-- -13
x"ffef0",-- -17
x"fff40",-- -12
x"fff40",-- -12
x"ffea0",-- -22
x"fff60",-- -10
x"00080",-- 8
x"00110",-- 17
x"00080",-- 8
x"fff40",-- -12
x"ffef0",-- -17
x"fff80",-- -8
x"00000",-- 0
x"000c0",-- 12
x"fff40",-- -12
x"ffe90",-- -23
x"fffb0",-- -5
x"fffb0",-- -5
x"fffe0",-- -2
x"fff80",-- -8
x"fff40",-- -12
x"ffec0",-- -20
x"fff80",-- -8
x"fffb0",-- -5
x"fffe0",-- -2
x"000c0",-- 12
x"fffb0",-- -5
x"fff40",-- -12
x"00020",-- 2
x"000f0",-- 15
x"00110",-- 17
x"000c0",-- 12
x"00140",-- 20
x"00170",-- 23
x"00160",-- 22
x"00120",-- 18
x"000c0",-- 12
x"00160",-- 22
x"001e0",-- 30
x"00200",-- 32
x"001e0",-- 30
x"001e0",-- 30
x"00210",-- 33
x"00140",-- 20
x"000c0",-- 12
x"000d0",-- 13
x"00020",-- 2
x"00020",-- 2
x"000a0",-- 10
x"00170",-- 23
x"00160",-- 22
x"00140",-- 20
x"000f0",-- 15
x"00020",-- 2
x"000f0",-- 15
x"00170",-- 23
x"001b0",-- 27
x"001e0",-- 30
x"00120",-- 18
x"00080",-- 8
x"00160",-- 22
x"00210",-- 33
x"001e0",-- 30
x"00160",-- 22
x"00160",-- 22
x"000a0",-- 10
x"000a0",-- 10
x"001e0",-- 30
x"00300",-- 48
x"00370",-- 55
x"002a0",-- 42
x"00250",-- 37
x"00230",-- 35
x"00300",-- 48
x"002a0",-- 42
x"00200",-- 32
x"00160",-- 22
x"000f0",-- 15
x"00190",-- 25
x"002b0",-- 43
x"002f0",-- 47
x"00230",-- 35
x"001c0",-- 28
x"001e0",-- 30
x"00250",-- 37
x"00300",-- 48
x"00280",-- 40
x"00230",-- 35
x"001e0",-- 30
x"00210",-- 33
x"00250",-- 37
x"001e0",-- 30
x"00210",-- 33
x"00170",-- 23
x"001c0",-- 28
x"00110",-- 17
x"00120",-- 18
x"001b0",-- 27
x"000f0",-- 15
x"00170",-- 23
x"00160",-- 22
x"00110",-- 17
x"000f0",-- 15
x"000c0",-- 12
x"00120",-- 18
x"000c0",-- 12
x"00080",-- 8
x"00050",-- 5
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00050",-- 5
x"000d0",-- 13
x"00050",-- 5
x"00020",-- 2
x"000a0",-- 10
x"00050",-- 5
x"000c0",-- 12
x"000a0",-- 10
x"00080",-- 8
x"000f0",-- 15
x"00120",-- 18
x"00140",-- 20
x"00160",-- 22
x"000f0",-- 15
x"00050",-- 5
x"00080",-- 8
x"000f0",-- 15
x"00160",-- 22
x"00120",-- 18
x"00110",-- 17
x"00120",-- 18
x"00160",-- 22
x"00050",-- 5
x"000f0",-- 15
x"001e0",-- 30
x"00080",-- 8
x"00160",-- 22
x"00070",-- 7
x"fffb0",-- -5
x"00000",-- 0
x"fffb0",-- -5
x"fff80",-- -8
x"fff40",-- -12
x"fff90",-- -7
x"fff80",-- -8
x"fff40",-- -12
x"ffef0",-- -17
x"fff10",-- -15
x"ffec0",-- -20
x"fff80",-- -8
x"ffef0",-- -17
x"fffe0",-- -2
x"00000",-- 0
x"fffd0",-- -3
x"fff80",-- -8
x"fff10",-- -15
x"fffb0",-- -5
x"fff80",-- -8
x"fffb0",-- -5
x"fff10",-- -15
x"fff10",-- -15
x"ffe00",-- -32
x"ffee0",-- -18
x"ffee0",-- -18
x"ffea0",-- -22
x"fff80",-- -8
x"ffe70",-- -25
x"ffee0",-- -18
x"ffe70",-- -25
x"ffea0",-- -22
x"ffdb0",-- -37
x"ffd50",-- -43
x"ffe20",-- -30
x"ffda0",-- -38
x"ffd80",-- -40
x"ffdb0",-- -37
x"ffd10",-- -47
x"ffc90",-- -55
x"ffc40",-- -60
x"ffc90",-- -55
x"ffd10",-- -47
x"ffda0",-- -38
x"ffdb0",-- -37
x"ffd10",-- -47
x"ffd60",-- -42
x"ffdb0",-- -37
x"ffdb0",-- -37
x"ffdb0",-- -37
x"ffd10",-- -47
x"ffd60",-- -42
x"ffd30",-- -45
x"ffd30",-- -45
x"ffdb0",-- -37
x"ffd30",-- -45
x"ffd30",-- -45
x"ffd30",-- -45
x"ffce0",-- -50
x"ffce0",-- -50
x"ffc90",-- -55
x"ffce0",-- -50
x"ffd10",-- -47
x"ffc10",-- -63
x"ffbc0",-- -68
x"ffb80",-- -72
x"ffc70",-- -57
x"ffce0",-- -50
x"ffc10",-- -63
x"ffbd0",-- -67
x"ffbf0",-- -65
x"ffbd0",-- -67
x"ffb20",-- -78
x"ffbc0",-- -68
x"ffb80",-- -72
x"ffbd0",-- -67
x"ffb50",-- -75
x"ffb20",-- -78
x"ffb50",-- -75
x"ffbf0",-- -65
x"ffb50",-- -75
x"ffbf0",-- -65
x"ffba0",-- -70
x"ffc60",-- -58
x"ffb50",-- -75
x"ffbd0",-- -67
x"ffef0",-- -17
x"ff940",-- -108
x"ffbf0",-- -65
x"ffd60",-- -42
x"ffc60",-- -58
x"ffda0",-- -38
x"ffcc0",-- -52
x"ffce0",-- -50
x"ffd50",-- -43
x"ffdb0",-- -37
x"ffce0",-- -50
x"ffd80",-- -40
x"ffda0",-- -38
x"ffd60",-- -42
x"ffdf0",-- -33
x"ffd50",-- -43
x"ffd10",-- -47
x"ffc90",-- -55
x"ffc90",-- -55
x"ffd10",-- -47
x"ffc60",-- -58
x"ffc10",-- -63
x"ffc20",-- -62
x"ffce0",-- -50
x"ffc90",-- -55
x"ffc90",-- -55
x"ffdb0",-- -37
x"ffd00",-- -48
x"ffc60",-- -58
x"ffd50",-- -43
x"ffda0",-- -38
x"ffdb0",-- -37
x"ffce0",-- -50
x"ffd30",-- -45
x"ffdf0",-- -33
x"ffdd0",-- -35
x"ffe20",-- -30
x"ffe00",-- -32
x"ffe50",-- -27
x"ffe50",-- -27
x"ffe40",-- -28
x"fff10",-- -15
x"fff60",-- -10
x"ffee0",-- -18
x"fff80",-- -8
x"00000",-- 0
x"00050",-- 5
x"00080",-- 8
x"00050",-- 5
x"00050",-- 5
x"00050",-- 5
x"000d0",-- 13
x"000c0",-- 12
x"000a0",-- 10
x"00110",-- 17
x"000c0",-- 12
x"000a0",-- 10
x"000d0",-- 13
x"00110",-- 17
x"000c0",-- 12
x"001b0",-- 27
x"00250",-- 37
x"002a0",-- 42
x"001b0",-- 27
x"00210",-- 33
x"002f0",-- 47
x"00250",-- 37
x"00280",-- 40
x"00210",-- 33
x"002a0",-- 42
x"001c0",-- 28
x"00210",-- 33
x"00280",-- 40
x"001e0",-- 30
x"001b0",-- 27
x"001e0",-- 30
x"00160",-- 22
x"00140",-- 20
x"000f0",-- 15
x"00080",-- 8
x"00020",-- 2
x"00000",-- 0
x"00000",-- 0
x"fff40",-- -12
x"fff90",-- -7
x"fff40",-- -12
x"fff40",-- -12
x"ffe20",-- -30
x"ffdf0",-- -33
x"ffdb0",-- -37
x"ffd60",-- -42
x"ffdf0",-- -33
x"ffd30",-- -45
x"ffd60",-- -42
x"ffd80",-- -40
x"ffdf0",-- -33
x"ffdd0",-- -35
x"ffe40",-- -28
x"ffdd0",-- -35
x"ffdf0",-- -33
x"ffe50",-- -27
x"ffea0",-- -22
x"ffee0",-- -18
x"ffe40",-- -28
x"ffea0",-- -22
x"ffe00",-- -32
x"ffe50",-- -27
x"ffec0",-- -20
x"ffee0",-- -18
x"ffea0",-- -22
x"ffda0",-- -38
x"ffdf0",-- -33
x"ffd30",-- -45
x"ffd80",-- -40
x"ffdf0",-- -33
x"ffce0",-- -50
x"ffc90",-- -55
x"ffcb0",-- -53
x"ffce0",-- -50
x"ffc70",-- -57
x"ffd30",-- -45
x"ffce0",-- -50
x"ffc90",-- -55
x"ffbf0",-- -65
x"ffb80",-- -72
x"ffc70",-- -57
x"ffbc0",-- -68
x"ffc20",-- -62
x"ffb80",-- -72
x"ffb20",-- -78
x"ffab0",-- -85
x"ffa60",-- -90
x"ffb00",-- -80
x"ffb20",-- -78
x"ffbd0",-- -67
x"ffb00",-- -80
x"ffab0",-- -85
x"ffa90",-- -87
x"ffa30",-- -93
x"ffad0",-- -83
x"ffa60",-- -90
x"ff9f0",-- -97
x"ff9e0",-- -98
x"ff9f0",-- -97
x"ffa60",-- -90
x"ff9f0",-- -97
x"ff950",-- -107
x"ff920",-- -110
x"ff9f0",-- -97
x"ff9a0",-- -102
x"ffad0",-- -83
x"ffa60",-- -90
x"ff9e0",-- -98
x"ffad0",-- -83
x"ffad0",-- -83
x"ffb20",-- -78
x"ffb00",-- -80
x"ffae0",-- -82
x"ffa90",-- -87
x"ffb20",-- -78
x"ffb50",-- -75
x"ffab0",-- -85
x"ffa60",-- -90
x"ffb00",-- -80
x"ffae0",-- -82
x"ffbc0",-- -68
x"ffb20",-- -78
x"ffb00",-- -80
x"ffb30",-- -77
x"ffa60",-- -90
x"ffb80",-- -72
x"ffb80",-- -72
x"ffb20",-- -78
x"ffae0",-- -82
x"ffa90",-- -87
x"ffb50",-- -75
x"ffa90",-- -87
x"ffad0",-- -83
x"ffb20",-- -78
x"ffa60",-- -90
x"ffa90",-- -87
x"ffad0",-- -83
x"ffb70",-- -73
x"ffb50",-- -75
x"ffb70",-- -73
x"ffae0",-- -82
x"ffb50",-- -75
x"ffa90",-- -87
x"ffb20",-- -78
x"ffc10",-- -63
x"ffc20",-- -62
x"ffce0",-- -50
x"ffcc0",-- -52
x"ffc90",-- -55
x"ffd10",-- -47
x"ffdf0",-- -33
x"ffdd0",-- -35
x"ffe70",-- -25
x"ffea0",-- -22
x"ffee0",-- -18
x"fff40",-- -12
x"fff40",-- -12
x"fff80",-- -8
x"00000",-- 0
x"fffd0",-- -3
x"fffe0",-- -2
x"00000",-- 0
x"fffe0",-- -2
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00160",-- 22
x"000a0",-- 10
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"000c0",-- 12
x"00070",-- 7
x"000f0",-- 15
x"00120",-- 18
x"00160",-- 22
x"00170",-- 23
x"00160",-- 22
x"001e0",-- 30
x"00160",-- 22
x"000f0",-- 15
x"00080",-- 8
x"000f0",-- 15
x"00250",-- 37
x"002b0",-- 43
x"001e0",-- 30
x"001c0",-- 28
x"00120",-- 18
x"000c0",-- 12
x"00140",-- 20
x"00160",-- 22
x"00120",-- 18
x"000c0",-- 12
x"00050",-- 5
x"00080",-- 8
x"00030",-- 3
x"00030",-- 3
x"000c0",-- 12
x"00050",-- 5
x"000c0",-- 12
x"00020",-- 2
x"000d0",-- 13
x"00170",-- 23
x"000f0",-- 15
x"000f0",-- 15
x"000c0",-- 12
x"000f0",-- 15
x"00120",-- 18
x"00230",-- 35
x"002b0",-- 43
x"00280",-- 40
x"00210",-- 33
x"00160",-- 22
x"001b0",-- 27
x"00250",-- 37
x"002a0",-- 42
x"00250",-- 37
x"002b0",-- 43
x"00250",-- 37
x"001e0",-- 30
x"001c0",-- 28
x"00110",-- 17
x"001b0",-- 27
x"00210",-- 33
x"00140",-- 20
x"00160",-- 22
x"00230",-- 35
x"001c0",-- 28
x"00210",-- 33
x"00200",-- 32
x"00250",-- 37
x"00210",-- 33
x"00160",-- 22
x"00210",-- 33
x"001e0",-- 30
x"001c0",-- 28
x"00210",-- 33
x"00210",-- 33
x"001e0",-- 30
x"00170",-- 23
x"001b0",-- 27
x"00160",-- 22
x"00230",-- 35
x"00210",-- 33
x"00190",-- 25
x"001e0",-- 30
x"001b0",-- 27
x"00280",-- 40
x"00280",-- 40
x"002b0",-- 43
x"00200",-- 32
x"00170",-- 23
x"00120",-- 18
x"00080",-- 8
x"00050",-- 5
x"00000",-- 0
x"00030",-- 3
x"000c0",-- 12
x"00050",-- 5
x"00050",-- 5
x"000d0",-- 13
x"000c0",-- 12
x"00120",-- 18
x"000f0",-- 15
x"00030",-- 3
x"00080",-- 8
x"000f0",-- 15
x"00140",-- 20
x"001b0",-- 27
x"000d0",-- 13
x"001e0",-- 30
x"00160",-- 22
x"001c0",-- 28
x"002a0",-- 42
x"001e0",-- 30
x"00230",-- 35
x"00260",-- 38
x"00210",-- 33
x"001b0",-- 27
x"00280",-- 40
x"002b0",-- 43
x"00300",-- 48
x"00280",-- 40
x"00210",-- 33
x"00210",-- 33
x"00230",-- 35
x"001e0",-- 30
x"001c0",-- 28
x"00210",-- 33
x"00280",-- 40
x"00200",-- 32
x"001c0",-- 28
x"00210",-- 33
x"00280",-- 40
x"00250",-- 37
x"001e0",-- 30
x"00280",-- 40
x"00210",-- 33
x"00200",-- 32
x"001e0",-- 30
x"001c0",-- 28
x"00210",-- 33
x"00210",-- 33
x"001e0",-- 30
x"001b0",-- 27
x"00160",-- 22
x"000a0",-- 10
x"000c0",-- 12
x"001b0",-- 27
x"00190",-- 25
x"000f0",-- 15
x"000f0",-- 15
x"000c0",-- 12
x"000c0",-- 12
x"00020",-- 2
x"000c0",-- 12
x"000f0",-- 15
x"000f0",-- 15
x"000f0",-- 15
x"001b0",-- 27
x"001b0",-- 27
x"00160",-- 22
x"000c0",-- 12
x"000d0",-- 13
x"001e0",-- 30
x"00110",-- 17
x"001b0",-- 27
x"00190",-- 25
x"00250",-- 37
x"00280",-- 40
x"001c0",-- 28
x"00250",-- 37
x"00280",-- 40
x"001b0",-- 27
x"001e0",-- 30
x"00120",-- 18
x"00140",-- 20
x"00200",-- 32
x"00110",-- 17
x"00070",-- 7
x"000f0",-- 15
x"00140",-- 20
x"000c0",-- 12
x"00080",-- 8
x"00030",-- 3
x"fffe0",-- -2
x"fff40",-- -12
x"fff30",-- -13
x"fff40",-- -12
x"fffb0",-- -5
x"ffee0",-- -18
x"ffe40",-- -28
x"ffdb0",-- -37
x"ffec0",-- -20
x"ffe40",-- -28
x"ffd80",-- -40
x"ffd80",-- -40
x"ffc70",-- -57
x"ffd30",-- -45
x"ffce0",-- -50
x"ffcb0",-- -53
x"ffc20",-- -62
x"ffc60",-- -58
x"ffc90",-- -55
x"ffc60",-- -58
x"ffcc0",-- -52
x"ffcc0",-- -52
x"ffd10",-- -47
x"ffd50",-- -43
x"ffdd0",-- -35
x"ffe20",-- -30
x"ffec0",-- -20
x"fff80",-- -8
x"00000",-- 0
x"00000",-- 0
x"fffe0",-- -2
x"000a0",-- 10
x"00000",-- 0
x"00020",-- 2
x"00080",-- 8
x"00080",-- 8
x"00120",-- 18
x"00160",-- 22
x"001c0",-- 28
x"00160",-- 22
x"000f0",-- 15
x"000c0",-- 12
x"000f0",-- 15
x"00080",-- 8
x"000c0",-- 12
x"00030",-- 3
x"00030",-- 3
x"000a0",-- 10
x"00000",-- 0
x"00020",-- 2
x"fff90",-- -7
x"ffe90",-- -23
x"ffea0",-- -22
x"ffe70",-- -25
x"ffd50",-- -43
x"ffc20",-- -62
x"ffb30",-- -77
x"ffb30",-- -77
x"ffa80",-- -88
x"ff9c0",-- -100
x"ff8d0",-- -115
x"ff710",-- -143
x"ff630",-- -157
x"ff600",-- -160
x"ff510",-- -175
x"ff4e0",-- -178
x"ff3b0",-- -197
x"ff350",-- -203
x"ff290",-- -215
x"ff260",-- -218
x"ff3a0",-- -198
x"ff380",-- -200
x"ff400",-- -192
x"ff470",-- -185
x"ff580",-- -168
x"ff6d0",-- -147
x"ff8b0",-- -117
x"ffa30",-- -93
x"ffb50",-- -75
x"ffc60",-- -58
x"ffe20",-- -30
x"00020",-- 2
x"00190",-- 25
x"003a0",-- 58
x"004e0",-- 78
x"00670",-- 103
x"00850",-- 133
x"00910",-- 145
x"00b20",-- 178
x"00c50",-- 197
x"00d90",-- 217
x"00e80",-- 232
x"00f20",-- 242
x"00fa0",-- 250
x"01080",-- 264
x"011a0",-- 282
x"011c0",-- 284
x"01220",-- 290
x"01260",-- 294
x"01100",-- 272
x"00d40",-- 212
x"00870",-- 135
x"00340",-- 52
x"00080",-- 8
x"00030",-- 3
x"fff10",-- -15
x"ffb20",-- -78
x"ff380",-- -200
x"fecb0",-- -309
x"fe840",-- -380
x"fe700",-- -400
x"fe580",-- -424
x"fe120",-- -494
x"fdc10",-- -575
x"fd6f0",-- -657
x"fd710",-- -655
x"fd9c0",-- -612
x"fdb50",-- -587
x"fda90",-- -599
x"fda40",-- -604
x"fdc20",-- -574
x"fe080",-- -504
x"fe710",-- -399
x"fed90",-- -295
x"ff330",-- -205
x"ff740",-- -140
x"ffce0",-- -50
x"002d0",-- 45
x"008f0",-- 143
x"00fa0",-- 250
x"015e0",-- 350
x"01a60",-- 422
x"01e50",-- 485
x"021c0",-- 540
x"02550",-- 597
x"02980",-- 664
x"02e00",-- 736
x"031a0",-- 794
x"03260",-- 806
x"032c0",-- 812
x"03400",-- 832
x"034c0",-- 844
x"034c0",-- 844
x"03540",-- 852
x"023e0",-- 574
x"003c0",-- 60
x"ff8a0",-- -118
x"00d50",-- 213
x"01e50",-- 485
x"00980",-- 152
x"fe890",-- -375
x"fd2e0",-- -722
x"fccf0",-- -817
x"fd850",-- -635
x"fe820",-- -382
x"fdda0",-- -550
x"fba40",-- -1116
x"fac30",-- -1341
x"fbc40",-- -1084
x"fcb90",-- -839
x"fd2c0",-- -724
x"fd9f0",-- -609
x"fd6c0",-- -660
x"fcfd0",-- -771
x"fddd0",-- -547
x"ff950",-- -107
x"00660",-- 102
x"00e40",-- 228
x"01c70",-- 455
x"021c0",-- 540
x"01db0",-- 475
x"02430",-- 579
x"03490",-- 841
x"03c60",-- 966
x"03ee0",-- 1006
x"03ce0",-- 974
x"02e30",-- 739
x"01ef0",-- 495
x"02120",-- 530
x"02870",-- 647
x"020f0",-- 527
x"010d0",-- 269
x"ffea0",-- -22
x"fec10",-- -319
x"fe2d0",-- -467
x"fe500",-- -432
x"fe3a0",-- -454
x"fd680",-- -664
x"fc820",-- -894
x"fbf80",-- -1032
x"fbc10",-- -1087
x"fbfd0",-- -1027
x"fc8f0",-- -881
x"fcdf0",-- -801
x"fcd40",-- -812
x"fcd70",-- -809
x"fd3a0",-- -710
x"fdcb0",-- -565
x"fea50",-- -347
x"ffa60",-- -90
x"00440",-- 68
x"00700",-- 112
x"00ac0",-- 172
x"01380",-- 312
x"01db0",-- 475
x"028e0",-- 654
x"03100",-- 784
x"03090",-- 777
x"02aa0",-- 682
x"02750",-- 629
x"02a00",-- 672
x"02d60",-- 726
x"02b10",-- 689
x"02500",-- 592
x"019a0",-- 410
x"00e30",-- 227
x"007b0",-- 123
x"00440",-- 68
x"000c0",-- 12
x"ff9f0",-- -97
x"ff170",-- -233
x"fe7a0",-- -390
x"fe0a0",-- -502
x"fdec0",-- -532
x"fdf60",-- -522
x"fe000",-- -512
x"fdf10",-- -527
x"fdd50",-- -555
x"fdc40",-- -572
x"fde70",-- -537
x"fe570",-- -425
x"fedf0",-- -289
x"ff440",-- -188
x"ff8a0",-- -118
x"ffad0",-- -83
x"ffe50",-- -27
x"00550",-- 85
x"00eb0",-- 235
x"01630",-- 355
x"01850",-- 389
x"01770",-- 375
x"01790",-- 377
x"018b0",-- 395
x"01c20",-- 450
x"01e40",-- 484
x"01cc0",-- 460
x"017b0",-- 379
x"011c0",-- 284
x"00d90",-- 217
x"00a80",-- 168
x"00850",-- 133
x"00530",-- 83
x"00000",-- 0
x"ff860",-- -122
x"ff270",-- -217
x"fef50",-- -267
x"feda0",-- -294
x"fec50",-- -315
x"feb40",-- -332
x"fe850",-- -379
x"fe5a0",-- -422
x"fe5d0",-- -419
x"fe760",-- -394
x"feb70",-- -329
x"fef70",-- -265
x"ff1f0",-- -225
x"ff3b0",-- -197
x"ff6a0",-- -150
x"ffb50",-- -75
x"00020",-- 2
x"00530",-- 83
x"00980",-- 152
x"00d50",-- 213
x"00f00",-- 240
x"01030",-- 259
x"012b0",-- 299
x"01510",-- 337
x"01630",-- 355
x"016a0",-- 362
x"01650",-- 357
x"013b0",-- 315
x"01130",-- 275
x"00f90",-- 249
x"00e80",-- 232
x"00d40",-- 212
x"00a30",-- 163
x"00460",-- 70
x"fffb0",-- -5
x"ffc70",-- -57
x"ffb00",-- -80
x"ffa60",-- -90
x"ff790",-- -135
x"ff3d0",-- -195
x"ff070",-- -249
x"fefd0",-- -259
x"ff010",-- -255
x"ff0e0",-- -242
x"ff110",-- -239
x"ff100",-- -240
x"ff0b0",-- -245
x"ff180",-- -232
x"ff4a0",-- -182
x"ff790",-- -135
x"ffad0",-- -83
x"ffd80",-- -40
x"ffee0",-- -18
x"000d0",-- 13
x"00440",-- 68
x"007a0",-- 122
x"00af0",-- 175
x"00dc0",-- 220
x"00e30",-- 227
x"00d70",-- 215
x"00e80",-- 232
x"00fc0",-- 252
x"00ff0",-- 255
x"00f90",-- 249
x"00dc0",-- 220
x"00b60",-- 182
x"00980",-- 152
x"00760",-- 118
x"00760",-- 118
x"00570",-- 87
x"00370",-- 55
x"000c0",-- 12
x"ffd80",-- -40
x"ffc10",-- -63
x"ffa80",-- -88
x"ff970",-- -105
x"ff790",-- -135
x"ff630",-- -157
x"ff510",-- -175
x"ff400",-- -192
x"ff470",-- -185
x"ff540",-- -172
x"ff560",-- -170
x"ff650",-- -155
x"ff7c0",-- -132
x"ff7c0",-- -132
x"ff950",-- -107
x"ffba0",-- -70
x"ffe50",-- -27
x"00050",-- 5
x"00120",-- 18
x"002b0",-- 43
x"00460",-- 70
x"00570",-- 87
x"008c0",-- 140
x"00aa0",-- 170
x"00ac0",-- 172
x"00a80",-- 168
x"00a80",-- 168
x"00940",-- 148
x"008e0",-- 142
x"00930",-- 147
x"007a0",-- 122
x"00530",-- 83
x"00300",-- 48
x"000d0",-- 13
x"ffec0",-- -20
x"ffd30",-- -45
x"ffc20",-- -62
x"ffad0",-- -83
x"ff940",-- -108
x"ff880",-- -120
x"ff720",-- -142
x"ff6d0",-- -147
x"ff6c0",-- -148
x"ff710",-- -143
x"ff6d0",-- -147
x"ff680",-- -152
x"ff790",-- -135
x"ff8d0",-- -115
x"ffb80",-- -72
x"ffda0",-- -38
x"fff10",-- -15
x"00000",-- 0
x"00160",-- 22
x"00370",-- 55
x"00480",-- 72
x"00530",-- 83
x"00730",-- 115
x"00820",-- 130
x"00800",-- 128
x"008f0",-- 143
x"00890",-- 137
x"008a0",-- 138
x"00850",-- 133
x"007b0",-- 123
x"00670",-- 103
x"00530",-- 83
x"004b0",-- 75
x"003a0",-- 58
x"00200",-- 32
x"00080",-- 8
x"fff90",-- -7
x"ffe20",-- -30
x"ffce0",-- -50
x"ffbd0",-- -67
x"ffb30",-- -77
x"ffb00",-- -80
x"ffa90",-- -87
x"ff990",-- -103
x"ff950",-- -107
x"ff9e0",-- -98
x"ffae0",-- -82
x"ffbf0",-- -65
x"ffc10",-- -63
x"ffcb0",-- -53
x"ffd80",-- -40
x"ffe40",-- -28
x"ffef0",-- -17
x"00000",-- 0
x"000c0",-- 12
x"000f0",-- 15
x"002b0",-- 43
x"002f0",-- 47
x"003a0",-- 58
x"00520",-- 82
x"00570",-- 87
x"006b0",-- 107
x"006e0",-- 110
x"00670",-- 103
x"00620",-- 98
x"00610",-- 97
x"00640",-- 100
x"00500",-- 80
x"00480",-- 72
x"00300",-- 48
x"00170",-- 23
x"00070",-- 7
x"fff90",-- -7
x"ffea0",-- -22
x"ffdf0",-- -33
x"ffd10",-- -47
x"ffc20",-- -62
x"ffb50",-- -75
x"ffa90",-- -87
x"ffb00",-- -80
x"ffae0",-- -82
x"ffad0",-- -83
x"ffb20",-- -78
x"ffb20",-- -78
x"ffc10",-- -63
x"ffcb0",-- -53
x"ffdb0",-- -37
x"ffee0",-- -18
x"ffe50",-- -27
x"fff30",-- -13
x"00030",-- 3
x"001b0",-- 27
x"00280",-- 40
x"00340",-- 52
x"00370",-- 55
x"00480",-- 72
x"00480",-- 72
x"00410",-- 65
x"00440",-- 68
x"00410",-- 65
x"00440",-- 68
x"00340",-- 52
x"002d0",-- 45
x"00210",-- 33
x"00120",-- 18
x"00050",-- 5
x"00000",-- 0
x"fff40",-- -12
x"ffdf0",-- -33
x"ffd10",-- -47
x"ffd10",-- -47
x"ffc20",-- -62
x"ffb20",-- -78
x"ffad0",-- -83
x"ffa30",-- -93
x"ffa60",-- -90
x"ffa40",-- -92
x"ffa80",-- -88
x"ffb50",-- -75
x"ffbc0",-- -68
x"ffcc0",-- -52
x"ffce0",-- -50
x"ffdd0",-- -35
x"ffee0",-- -18
x"00000",-- 0
x"00000",-- 0
x"00080",-- 8
x"00250",-- 37
x"00210",-- 33
x"00340",-- 52
x"00410",-- 65
x"004b0",-- 75
x"00500",-- 80
x"004b0",-- 75
x"00410",-- 65
x"00320",-- 50
x"002b0",-- 43
x"00370",-- 55
x"00250",-- 37
x"00140",-- 20
x"00000",-- 0
x"fff10",-- -15
x"fff80",-- -8
x"ffe20",-- -30
x"ffd30",-- -45
x"ffc90",-- -55
x"ffbf0",-- -65
x"ffc40",-- -60
x"ffc40",-- -60
x"ffc90",-- -55
x"ffc90",-- -55
x"ffc60",-- -58
x"ffc20",-- -62
x"ffc20",-- -62
x"ffd50",-- -43
x"ffe40",-- -28
x"fff60",-- -10
x"00030",-- 3
x"00050",-- 5
x"00050",-- 5
x"000f0",-- 15
x"00210",-- 33
x"00250",-- 37
x"002b0",-- 43
x"002f0",-- 47
x"00320",-- 50
x"00350",-- 53
x"002f0",-- 47
x"00350",-- 53
x"00370",-- 55
x"00370",-- 55
x"00340",-- 52
x"00250",-- 37
x"001e0",-- 30
x"00110",-- 17
x"00080",-- 8
x"00070",-- 7
x"fffb0",-- -5
x"ffee0",-- -18
x"ffea0",-- -22
x"ffe90",-- -23
x"ffe50",-- -27
x"ffea0",-- -22
x"ffe20",-- -30
x"ffdb0",-- -37
x"ffe20",-- -30
x"ffd80",-- -40
x"ffe50",-- -27
x"ffe20",-- -30
x"ffe00",-- -32
x"ffe90",-- -23
x"ffee0",-- -18
x"fffb0",-- -5
x"00000",-- 0
x"00070",-- 7
x"00050",-- 5
x"000c0",-- 12
x"000f0",-- 15
x"00200",-- 32
x"002b0",-- 43
x"00280",-- 40
x"00280",-- 40
x"002b0",-- 43
x"003a0",-- 58
x"003e0",-- 62
x"00340",-- 52
x"002b0",-- 43
x"00210",-- 33
x"00250",-- 37
x"00250",-- 37
x"00210",-- 33
x"00080",-- 8
x"00020",-- 2
x"000d0",-- 13
x"00070",-- 7
x"00020",-- 2
x"fffb0",-- -5
x"fff40",-- -12
x"ffec0",-- -20
x"ffea0",-- -22
x"ffef0",-- -17
x"fff40",-- -12
x"ffef0",-- -17
x"fff10",-- -15
x"fff60",-- -10
x"fff40",-- -12
x"fffe0",-- -2
x"fffb0",-- -5
x"00000",-- 0
x"00000",-- 0
x"fffd0",-- -3
x"00000",-- 0
x"00000",-- 0
x"000c0",-- 12
x"00110",-- 17
x"00160",-- 22
x"00200",-- 32
x"00190",-- 25
x"00120",-- 18
x"001b0",-- 27
x"000c0",-- 12
x"000c0",-- 12
x"000c0",-- 12
x"00000",-- 0
x"fff60",-- -10
x"ffef0",-- -17
x"fff30",-- -13
x"ffef0",-- -17
x"fff10",-- -15
x"ffe70",-- -25
x"ffd50",-- -43
x"ffd10",-- -47
x"ffd60",-- -42
x"ffd00",-- -48
x"ffd10",-- -47
x"ffcb0",-- -53
x"ffcb0",-- -53
x"ffcc0",-- -52
x"ffc40",-- -60
x"ffcb0",-- -53
x"ffc70",-- -57
x"ffc90",-- -55
x"ffcc0",-- -52
x"ffcc0",-- -52
x"ffd60",-- -42
x"ffe20",-- -30
x"ffe50",-- -27
x"ffe90",-- -23
x"ffe70",-- -25
x"ffea0",-- -22
x"ffef0",-- -17
x"fff40",-- -12
x"fff30",-- -13
x"fff80",-- -8
x"fffb0",-- -5
x"fff30",-- -13
x"fff10",-- -15
x"fff60",-- -10
x"fff40",-- -12
x"ffef0",-- -17
x"fff40",-- -12
x"ffef0",-- -17
x"ffee0",-- -18
x"ffea0",-- -22
x"ffea0",-- -22
x"ffdb0",-- -37
x"ffdf0",-- -33
x"ffe40",-- -28
x"ffd60",-- -42
x"ffdf0",-- -33
x"ffdf0",-- -33
x"fff10",-- -15
x"ffee0",-- -18
x"fff10",-- -15
x"fff10",-- -15
x"ffee0",-- -18
x"fff80",-- -8
x"00000",-- 0
x"00020",-- 2
x"00050",-- 5
x"00000",-- 0
x"fffb0",-- -5
x"fff90",-- -7
x"fff80",-- -8
x"00000",-- 0
x"00000",-- 0
x"000f0",-- 15
x"00080",-- 8
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fffe0",-- -2
x"00020",-- 2
x"00050",-- 5
x"fff90",-- -7
x"00070",-- 7
x"fffe0",-- -2
x"fffd0",-- -3
x"fffd0",-- -3
x"fffe0",-- -2
x"fffe0",-- -2
x"fffe0",-- -2
x"00020",-- 2
x"00080",-- 8
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fffe0",-- -2
x"00030",-- 3
x"00000",-- 0
x"00030",-- 3
x"fffb0",-- -5
x"00000",-- 0
x"fffb0",-- -5
x"fffb0",-- -5
x"00000",-- 0
x"fffb0",-- -5
x"00050",-- 5
x"00050",-- 5
x"00030",-- 3
x"fff60",-- -10
x"fffe0",-- -2
x"ffef0",-- -17
x"00110",-- 17
x"ffe00",-- -32
x"ff8b0",-- -117
x"ffe20",-- -30
x"fffd0",-- -3
x"00000",-- 0
x"ffbc0",-- -68
x"ff8a0",-- -118
x"ff6a0",-- -150
x"ff8b0",-- -117
x"ffce0",-- -50
x"ffa10",-- -95
x"ff150",-- -235
x"fec30",-- -317
x"ff220",-- -222
x"ff970",-- -105
x"ff6a0",-- -150
x"fef00",-- -272
x"fe9e0",-- -354
x"fe8c0",-- -372
x"fe840",-- -380
x"fe340",-- -460
x"fe3f0",-- -449
x"fdae0",-- -594
x"fdf60",-- -522
x"fe340",-- -460
x"fe2a0",-- -470
x"fdc10",-- -575
x"fd680",-- -664
x"fdfb0",-- -517
x"fe460",-- -442
x"feaf0",-- -337
x"fe530",-- -429
x"fe1b0",-- -485
x"fe7a0",-- -390
x"ff240",-- -220
x"000d0",-- 13
x"00370",-- 55
x"ffd30",-- -45
x"00230",-- 35
x"00870",-- 135
x"01810",-- 385
x"01fe0",-- 510
x"02550",-- 597
x"02640",-- 612
x"025f0",-- 607
x"035e0",-- 862
x"03920",-- 914
x"042a0",-- 1066
x"04140",-- 1044
x"04710",-- 1137
x"04f90",-- 1273
x"057e0",-- 1406
x"06250",-- 1573
x"06d70",-- 1751
x"076a0",-- 1898
x"08550",-- 2133
x"08610",-- 2145
x"085e0",-- 2142
x"08c00",-- 2240
x"099c0",-- 2460
x"09f30",-- 2547
x"095b0",-- 2395
x"09090",-- 2313
x"05d00",-- 1488
x"04d60",-- 1238
x"04f40",-- 1268
x"06210",-- 1569
x"04550",-- 1109
x"00ef0",-- 239
x"fe930",-- -365
x"fc490",-- -951
x"fc4d0",-- -947
x"fbe90",-- -1047
x"fac50",-- -1339
x"f7950",-- -2155
x"f5540",-- -2732
x"f5010",-- -2815
x"f52e0",-- -2770
x"f57e0",-- -2690
x"f6300",-- -2512
x"f61e0",-- -2530
x"f6200",-- -2528
x"f6cf0",-- -2353
x"f8aa0",-- -1878
x"fa960",-- -1386
x"fc260",-- -986
x"fe460",-- -442
x"ffa60",-- -90
x"00d50",-- 213
x"017e0",-- 382
x"03290",-- 809
x"04a50",-- 1189
x"05c20",-- 1474
x"067f0",-- 1663
x"06610",-- 1633
x"057c0",-- 1404
x"04bb0",-- 1211
x"04fc0",-- 1276
x"04c70",-- 1223
x"03bc0",-- 956
x"02390",-- 569
x"00760",-- 118
x"fe710",-- -399
x"fd340",-- -716
x"fc9e0",-- -866
x"fba30",-- -1117
x"f9fe0",-- -1538
x"f8c50",-- -1851
x"f7660",-- -2202
x"f6480",-- -2488
x"f6570",-- -2473
x"f7100",-- -2288
x"f7510",-- -2223
x"f6f00",-- -2320
x"f6d70",-- -2345
x"f75c0",-- -2212
x"f8c10",-- -1855
x"fafc0",-- -1284
x"fc820",-- -894
x"fd160",-- -746
x"fdb20",-- -590
x"ff0c0",-- -244
x"009b0",-- 155
x"01ee0",-- 494
x"03da0",-- 986
x"04ae0",-- 1198
x"04ed0",-- 1261
x"050d0",-- 1293
x"05880",-- 1416
x"06260",-- 1574
x"062d0",-- 1581
x"06350",-- 1589
x"056c0",-- 1388
x"04440",-- 1092
x"035d0",-- 861
x"02f40",-- 756
x"027f0",-- 639
x"01830",-- 387
x"006c0",-- 108
x"ff2c0",-- -212
x"fdee0",-- -530
x"fd4c0",-- -692
x"fcf30",-- -781
x"fc690",-- -919
x"fbb70",-- -1097
x"fb570",-- -1193
x"fb5e0",-- -1186
x"fb680",-- -1176
x"fba60",-- -1114
x"fc000",-- -1024
x"fc750",-- -907
x"fd400",-- -704
x"fe140",-- -492
x"feb10",-- -335
x"ff440",-- -188
x"ffe90",-- -23
x"01030",-- 259
x"01bf0",-- 447
x"026b0",-- 619
x"02d60",-- 726
x"02e60",-- 742
x"031c0",-- 796
x"03760",-- 886
x"03fb0",-- 1019
x"03e50",-- 997
x"03330",-- 819
x"02aa0",-- 682
x"02350",-- 565
x"02280",-- 552
x"01bf0",-- 447
x"01210",-- 289
x"00530",-- 83
x"ff830",-- -125
x"ff380",-- -200
x"fe760",-- -394
x"fe480",-- -440
x"fde40",-- -540
x"fdd80",-- -552
x"fdad0",-- -595
x"fd060",-- -762
x"fd590",-- -679
x"fd530",-- -685
x"fe000",-- -512
x"fe1b0",-- -485
x"fe850",-- -379
x"feeb0",-- -277
x"ff4c0",-- -180
x"00700",-- 112
x"00640",-- 100
x"01180",-- 280
x"01950",-- 405
x"01db0",-- 475
x"024d0",-- 589
x"02ea0",-- 746
x"035b0",-- 859
x"02fa0",-- 762
x"034e0",-- 846
x"03ae0",-- 942
x"03bd0",-- 957
x"03f80",-- 1016
x"03830",-- 899
x"03850",-- 901
x"03130",-- 787
x"03210",-- 801
x"036a0",-- 874
x"03090",-- 777
x"034f0",-- 847
x"01d00",-- 464
x"02bc0",-- 700
x"03290",-- 809
x"03420",-- 834
x"03880",-- 904
x"03a10",-- 929
x"049b0",-- 1179
x"04e10",-- 1249
x"06b90",-- 1721
x"07850",-- 1925
x"079c0",-- 1948
x"06fa0",-- 1786
x"08b60",-- 2230
x"098d0",-- 2445
x"0c1e0",-- 3102
x"0d2c0",-- 3372
x"0e750",-- 3701
x"0b580",-- 2904
x"04300",-- 1072
x"03f90",-- 1017
x"05d60",-- 1494
x"0afa0",-- 2810
x"07ba0",-- 1978
x"01510",-- 337
x"fb380",-- -1224
x"f8550",-- -1963
x"fa620",-- -1438
x"fbc70",-- -1081
x"fa160",-- -1514
x"f36d0",-- -3219
x"eeda0",-- -4390
x"eed90",-- -4391
x"f10b0",-- -3829
x"f2280",-- -3544
x"f25c0",-- -3492
x"f0ee0",-- -3858
x"f1100",-- -3824
x"f2d90",-- -3367
x"f6250",-- -2523
x"f8410",-- -1983
x"f9a40",-- -1628
x"fc940",-- -876
x"febb0",-- -325
x"00d40",-- 212
x"01830",-- 387
x"028a0",-- 650
x"030d0",-- 781
x"04c30",-- 1219
x"06960",-- 1686
x"06020",-- 1538
x"039a0",-- 922
x"01a90",-- 425
x"00df0",-- 223
x"00c80",-- 200
x"00500",-- 80
x"fe460",-- -442
x"fa980",-- -1384
x"f74a0",-- -2230
x"f6000",-- -2560
x"f5da0",-- -2598
x"f52c0",-- -2772
x"f3900",-- -3184
x"f2050",-- -3579
x"f0eb0",-- -3861
x"f0fa0",-- -3846
x"f1f60",-- -3594
x"f3420",-- -3262
x"f4140",-- -3052
x"f5570",-- -2729
x"f7430",-- -2237
x"f92c0",-- -1748
x"fad20",-- -1326
x"fcda0",-- -806
x"ff0e0",-- -242
x"01b70",-- 439
x"04080",-- 1032
x"05ce0",-- 1486
x"07310",-- 1841
x"07d50",-- 2005
x"09ad0",-- 2477
x"0b4f0",-- 2895
x"0cd90",-- 3289
x"0d270",-- 3367
x"0d620",-- 3426
x"0dd10",-- 3537
x"0e7c0",-- 3708
x"0fa10",-- 4001
x"107c0",-- 4220
x"10750",-- 4213
x"0ff50",-- 4085
x"10d20",-- 4306
x"119c0",-- 4508
x"13770",-- 4983
x"13920",-- 5010
x"14b60",-- 5302
x"118a0",-- 4490
x"0ed40",-- 3796
x"0f650",-- 3941
x"0d220",-- 3362
x"0aea0",-- 2794
x"03bf0",-- 959
x"00490",-- 73
x"001b0",-- 27
x"00700",-- 112
x"fea70",-- -345
x"f75b0",-- -2213
x"f04e0",-- -4018
x"ebce0",-- -5170
x"ec740",-- -5004
x"ee640",-- -4508
x"ed150",-- -4843
x"e9040",-- -5884
x"e5ea0",-- -6678
x"e6c90",-- -6455
x"eb200",-- -5344
x"ef270",-- -4313
x"f1bf0",-- -3649
x"f3010",-- -3327
x"f4ff0",-- -2817
x"fa070",-- -1529
x"ff830",-- -125
x"03a80",-- 936
x"061e0",-- 1566
x"08d60",-- 2262
x"0b970",-- 2967
x"0e7c0",-- 3708
x"0f6d0",-- 3949
x"0ee80",-- 3816
x"0dd80",-- 3544
x"0da30",-- 3491
x"0d970",-- 3479
x"0b4f0",-- 2895
x"06760",-- 1654
x"02200",-- 544
x"00260",-- 38
x"fdb80",-- -584
x"fb3b0",-- -1221
x"f6490",-- -2487
x"f16d0",-- -3731
x"eda20",-- -4702
x"ebe30",-- -5149
x"ec420",-- -5054
x"eb2f0",-- -5329
x"e9330",-- -5837
x"e7630",-- -6301
x"e81c0",-- -6116
x"eadc0",-- -5412
x"ee380",-- -4552
x"f0c00",-- -3904
x"f25f0",-- -3489
x"f4730",-- -2957
x"f8eb0",-- -1813
x"fd900",-- -624
x"01b80",-- 440
x"04780",-- 1144
x"06820",-- 1666
x"09ad0",-- 2477
x"0c610",-- 3169
x"0efc0",-- 3836
x"0fb50",-- 4021
x"0fb80",-- 4024
x"0f490",-- 3913
x"0fd50",-- 4053
x"0f4c0",-- 3916
x"0df30",-- 3571
x"0bce0",-- 3022
x"09490",-- 2377
x"07ae0",-- 1966
x"05b80",-- 1464
x"042b0",-- 1067
x"01290",-- 297
x"ff2c0",-- -212
x"fd590",-- -679
x"fd160",-- -746
x"fcdf0",-- -801
x"fc530",-- -941
x"fcc60",-- -826
x"fd9f0",-- -609
x"ff270",-- -217
x"015e0",-- 350
x"05310",-- 1329
x"06fe0",-- 1790
x"0b0e0",-- 2830
x"0d830",-- 3459
x"10dc0",-- 4316
x"13e60",-- 5094
x"17490",-- 5961
x"1aa40",-- 6820
x"1d3a0",-- 7482
x"1eea0",-- 7914
x"22d40",-- 8916
x"1de70",-- 7655
x"0ce30",-- 3299
x"07240",-- 1828
x"0cbd0",-- 3261
x"162f0",-- 5679
x"12230",-- 4643
x"05580",-- 1368
x"f6850",-- -2427
x"ea230",-- -5597
x"eae10",-- -5407
x"f1ea0",-- -3606
x"f1f20",-- -3598
x"e5840",-- -6780
x"dadc0",-- -9508
x"d98b0",-- -9845
x"dd0a0",-- -8950
x"e16a0",-- -7830
x"e5860",-- -6778
x"e4b20",-- -6990
x"e3f20",-- -7182
x"ea0f0",-- -5617
x"f2c50",-- -3387
x"f8580",-- -1960
x"f9fe0",-- -1538
x"fe490",-- -439
x"041e0",-- 1054
x"0a1c0",-- 2588
x"0e0a0",-- 3594
x"10a50",-- 4261
x"0eff0",-- 3839
x"0e3b0",-- 3643
x"115e0",-- 4446
x"12cf0",-- 4815
x"11010",-- 4353
x"0c630",-- 3171
x"06dc0",-- 1756
x"02910",-- 657
x"fffe0",-- -2
x"feda0",-- -294
x"faca0",-- -1334
x"f39a0",-- -3174
x"eee60",-- -4378
x"ec1f0",-- -5089
x"ea6a0",-- -5526
x"e8da0",-- -5926
x"e7c00",-- -6208
x"e6300",-- -6608
x"e59c0",-- -6756
x"e8490",-- -6071
x"eb4c0",-- -5300
x"ec620",-- -5022
x"ee530",-- -4525
x"f2370",-- -3529
x"f7100",-- -2288
x"fc760",-- -906
x"00a80",-- 168
x"035d0",-- 861
x"04b40",-- 1204
x"08640",-- 2148
x"0db00",-- 3504
x"11100",-- 4368
x"11c10",-- 4545
x"117b0",-- 4475
x"10b80",-- 4280
x"10960",-- 4246
x"11940",-- 4500
x"11dc0",-- 4572
x"10b60",-- 4278
x"0e870",-- 3719
x"0dc70",-- 3527
x"0d240",-- 3364
x"0c480",-- 3144
x"0bd10",-- 3025
x"0b6f0",-- 2927
x"0c820",-- 3202
x"0df30",-- 3571
x"0f1a0",-- 3866
x"0f9a0",-- 3994
x"104b0",-- 4171
x"11c90",-- 4553
x"15800",-- 5504
x"18ed0",-- 6381
x"18050",-- 6149
x"16f50",-- 5877
x"12f90",-- 4857
x"0fd20",-- 4050
x"0ddd0",-- 3549
x"0a6e0",-- 2670
x"08d70",-- 2263
x"05450",-- 1349
x"01cc0",-- 460
x"fd6f0",-- -657
x"f6ca0",-- -2358
x"efd10",-- -4143
x"e8f80",-- -5896
x"e6be0",-- -6466
x"e5720",-- -6798
x"e4410",-- -7103
x"e1c90",-- -7735
x"def50",-- -8459
x"de1a0",-- -8678
x"e0800",-- -8064
x"e4c80",-- -6968
x"e8e90",-- -5911
x"ec600",-- -5024
x"f00b0",-- -4085
x"f56a0",-- -2710
x"fae30",-- -1309
x"00da0",-- 218
x"06460",-- 1606
x"0a370",-- 2615
x"0d810",-- 3457
x"0f740",-- 3956
x"0e540",-- 3668
x"0d6c0",-- 3436
x"0f790",-- 3961
x"11400",-- 4416
x"10680",-- 4200
x"0b6d0",-- 2925
x"062b0",-- 1579
x"00eb0",-- 235
x"fdab0",-- -597
x"fbb30",-- -1101
x"f78d0",-- -2163
x"f1a70",-- -3673
x"ec670",-- -5017
x"e9600",-- -5792
x"e71b0",-- -6373
x"e56b0",-- -6805
x"e39d0",-- -7267
x"e2960",-- -7530
x"e20f0",-- -7665
x"e4a60",-- -7002
x"e8280",-- -6104
x"ea460",-- -5562
x"ecd70",-- -4905
x"f0260",-- -4058
x"f5750",-- -2699
x"fa460",-- -1466
x"ff180",-- -232
x"03180",-- 792
x"06370",-- 1591
x"09470",-- 2375
x"0d650",-- 3429
x"10660",-- 4198
x"12780",-- 4728
x"13910",-- 5009
x"13ba0",-- 5050
x"141d0",-- 5149
x"12eb0",-- 4843
x"12400",-- 4672
x"100f0",-- 4111
x"0e0f0",-- 3599
x"0cd40",-- 3284
x"0c4a0",-- 3146
x"0afe0",-- 2814
x"08b30",-- 2227
x"07600",-- 1888
x"05bd0",-- 1469
x"05e50",-- 1509
x"07a30",-- 1955
x"0a520",-- 2642
x"0b940",-- 2964
x"0ce80",-- 3304
x"0ea20",-- 3746
x"11290",-- 4393
x"14dc0",-- 5340
x"19320",-- 6450
x"1c140",-- 7188
x"1acd0",-- 6861
x"1ba00",-- 7072
x"18480",-- 6216
x"155f0",-- 5471
x"11fd0",-- 4605
x"0ea50",-- 3749
x"0bf10",-- 3057
x"07c60",-- 1990
x"05d10",-- 1489
x"ff9a0",-- -102
x"f7750",-- -2187
x"ef3b0",-- -4293
x"ea910",-- -5487
x"e7020",-- -6398
x"e4ba0",-- -6982
x"e2c60",-- -7482
x"df6d0",-- -8339
x"dc580",-- -9128
x"dbb60",-- -9290
x"df140",-- -8428
x"e1a20",-- -7774
x"e5d10",-- -6703
x"e9880",-- -5752
x"ee550",-- -4523
x"f3510",-- -3247
x"f8c80",-- -1848
x"ff070",-- -249
x"03490",-- 841
x"075b0",-- 1883
x"09b00",-- 2480
x"0bcb0",-- 3019
x"0ec70",-- 3783
x"11e70",-- 4583
x"12310",-- 4657
x"105f0",-- 4191
x"0ceb0",-- 3307
x"0aa70",-- 2727
x"093d0",-- 2365
x"063a0",-- 1594
x"02280",-- 552
x"fb970",-- -1129
x"f62b0",-- -2517
x"f2520",-- -3502
x"ef310",-- -4303
x"ec3f0",-- -5057
x"e7e00",-- -6176
x"e4870",-- -7033
x"e2aa0",-- -7510
x"e2eb0",-- -7445
x"e4100",-- -7152
x"e5520",-- -6830
x"e66c0",-- -6548
x"e8a80",-- -5976
x"ecd50",-- -4907
x"f18b0",-- -3701
x"f5f60",-- -2570
x"f9590",-- -1703
x"fd6c0",-- -660
x"01db0",-- 475
x"06890",-- 1673
x"0b240",-- 2852
x"0dd60",-- 3542
x"0fc80",-- 4040
x"11bf0",-- 4543
x"13e20",-- 5090
x"151f0",-- 5407
x"15270",-- 5415
x"14390",-- 5177
x"12bd0",-- 4797
x"11620",-- 4450
x"107c0",-- 4220
x"0f9c0",-- 3996
x"0e460",-- 3654
x"0ca40",-- 3236
x"0b990",-- 2969
x"09c20",-- 2498
x"0a360",-- 2614
x"0b880",-- 2952
x"0d800",-- 3456
x"0db30",-- 3507
x"0e7d0",-- 3709
x"10bd0",-- 4285
x"12390",-- 4665
x"17940",-- 6036
x"19790",-- 6521
x"1a960",-- 6806
x"1a4d0",-- 6733
x"1da60",-- 7590
x"20640",-- 8292
x"1b320",-- 6962
x"146b0",-- 5227
x"0ea70",-- 3751
x"0b850",-- 2949
x"09510",-- 2385
x"089b0",-- 2203
x"05210",-- 1313
x"fbf60",-- -1034
x"f14a0",-- -3766
x"ebb00",-- -5200
x"e7b10",-- -6223
x"e3c40",-- -7228
x"e0a50",-- -8027
x"dd6b0",-- -8853
x"db250",-- -9435
x"d9a50",-- -9819
x"dbea0",-- -9238
x"dd190",-- -8935
x"dd750",-- -8843
x"e0fb0",-- -7941
x"e77e0",-- -6274
x"ee6b0",-- -4501
x"f47f0",-- -2945
x"fa0f0",-- -1521
x"fdab0",-- -597
x"00be0",-- 190
x"043f0",-- 1087
x"09740",-- 2420
x"0e200",-- 3616
x"11680",-- 4456
x"12870",-- 4743
x"10930",-- 4243
x"0de50",-- 3557
x"0bfd0",-- 3069
x"0aed0",-- 2797
x"07ef0",-- 2031
x"04340",-- 1076
x"ffbc0",-- -68
x"fa840",-- -1404
x"f5750",-- -2699
x"f0ff0",-- -3841
x"ecf50",-- -4875
x"e8cd0",-- -5939
x"e5cf0",-- -6705
x"e47b0",-- -7045
x"e3520",-- -7342
x"e1b30",-- -7757
x"e1ac0",-- -7764
x"e2a30",-- -7517
x"e4f30",-- -6925
x"e8f20",-- -5902
x"ed3d0",-- -4803
x"f0820",-- -3966
x"f4160",-- -3050
x"f8c60",-- -1850
x"fd880",-- -632
x"01f60",-- 502
x"069f0",-- 1695
x"0aa70",-- 2727
x"0e2c0",-- 3628
x"119e0",-- 4510
x"13e40",-- 5092
x"15830",-- 5507
x"15580",-- 5464
x"15bf0",-- 5567
x"15f50",-- 5621
x"157d0",-- 5501
x"15420",-- 5442
x"13920",-- 5010
x"11860",-- 4486
x"0fc40",-- 4036
x"0df30",-- 3571
x"0c9b0",-- 3227
x"0ca40",-- 3236
x"0df00",-- 3568
x"0e680",-- 3688
x"0e4d0",-- 3661
x"0e980",-- 3736
x"0e730",-- 3699
x"10590",-- 4185
x"13560",-- 4950
x"17370",-- 5943
x"1af10",-- 6897
x"1c070",-- 7175
x"1b0f0",-- 6927
x"1dd30",-- 7635
x"1e7f0",-- 7807
x"1ccf0",-- 7375
x"16780",-- 5752
x"11130",-- 4371
x"0d810",-- 3457
x"09bd0",-- 2493
x"08c00",-- 2240
x"06080",-- 1544
x"fe9b0",-- -357
x"f4260",-- -3034
x"ee850",-- -4475
x"e9220",-- -5854
x"e4f30",-- -6925
x"e11b0",-- -7909
x"de210",-- -8671
x"db2d0",-- -9427
x"d8c30",-- -10045
x"db720",-- -9358
x"dbcf0",-- -9265
x"dc530",-- -9133
x"de1a0",-- -8678
x"e3110",-- -7407
x"e8be0",-- -5954
x"eeb60",-- -4426
x"f54d0",-- -2739
x"f90b0",-- -1781
x"fa190",-- -1511
x"fe670",-- -409
x"05860",-- 1414
x"09ce0",-- 2510
x"0d760",-- 3446
x"0dfd0",-- 3581
x"0d8a0",-- 3466
x"0c640",-- 3172
x"0c270",-- 3111
x"0bf60",-- 3062
x"08440",-- 2116
x"04230",-- 1059
x"022f0",-- 559
x"fef50",-- -267
x"fb090",-- -1271
x"f6c60",-- -2362
x"f17f0",-- -3713
x"ecbc0",-- -4932
x"e97e0",-- -5762
x"e93b0",-- -5829
x"e7dd0",-- -6179
x"e5880",-- -6776
x"e4880",-- -7032
x"e4d00",-- -6960
x"e5a20",-- -6750
x"e8a10",-- -5983
x"ebf70",-- -5129
x"eeaa0",-- -4438
x"f1a70",-- -3673
x"f5f30",-- -2573
x"fadc0",-- -1316
x"fdef0",-- -529
x"021b0",-- 539
x"06050",-- 1541
x"096f0",-- 2415
x"0dda0",-- 3546
x"10f00",-- 4336
x"12e30",-- 4835
x"130d0",-- 4877
x"13710",-- 4977
x"14750",-- 5237
x"15670",-- 5479
x"16360",-- 5686
x"162c0",-- 5676
x"14cf0",-- 5327
x"12f40",-- 4852
x"11e10",-- 4577
x"11030",-- 4355
x"10b90",-- 4281
x"11a60",-- 4518
x"122d0",-- 4653
x"117e0",-- 4478
x"11180",-- 4376
x"110d0",-- 4365
x"12e30",-- 4835
x"14b10",-- 5297
x"182a0",-- 6186
x"1b210",-- 6945
x"1b920",-- 7058
x"1b080",-- 6920
x"1ad60",-- 6870
x"1c610",-- 7265
x"1c500",-- 7248
x"17e70",-- 6119
x"13090",-- 4873
x"0f590",-- 3929
x"0cb10",-- 3249
x"09760",-- 2422
x"059f0",-- 1439
x"00840",-- 132
x"f92a0",-- -1750
x"f3e50",-- -3099
x"efbb0",-- -4165
x"ea9c0",-- -5476
x"e4c30",-- -6973
x"e0260",-- -8154
x"dda00",-- -8800
x"db6e0",-- -9362
x"db910",-- -9327
x"dc460",-- -9146
x"dc1f0",-- -9185
x"dc060",-- -9210
x"df430",-- -8381
x"e3890",-- -7287
x"e7ab0",-- -6229
x"eb810",-- -5247
x"eeff0",-- -4353
x"f38e0",-- -3186
x"f8990",-- -1895
x"fe820",-- -382
x"02030",-- 515
x"03850",-- 901
x"051f0",-- 1311
x"076d0",-- 1901
x"09170",-- 2327
x"0a700",-- 2672
x"09e00",-- 2528
x"07580",-- 1880
x"05240",-- 1316
x"03b50",-- 949
x"02f50",-- 757
x"ffdb0",-- -37
x"fbe00",-- -1056
x"f7f10",-- -2063
x"f45a0",-- -2982
x"f21c0",-- -3556
x"f0190",-- -4071
x"eda70",-- -4697
x"ea620",-- -5534
x"e95c0",-- -5796
x"e97a0",-- -5766
x"ea620",-- -5534
x"eabe0",-- -5442
x"eba90",-- -5207
x"ecb60",-- -4938
x"ee710",-- -4495
x"f2a20",-- -3422
x"f5fe0",-- -2562
x"f9680",-- -1688
x"fbf80",-- -1032
x"ffc10",-- -63
x"036f0",-- 879
x"07170",-- 1815
x"0ab40",-- 2740
x"0cf90",-- 3321
x"0f150",-- 3861
x"11450",-- 4421
x"13ba0",-- 5050
x"153b0",-- 5435
x"16550",-- 5717
x"167d0",-- 5757
x"169b0",-- 5787
x"16570",-- 5719
x"160f0",-- 5647
x"15920",-- 5522
x"14e00",-- 5344
x"14570",-- 5207
x"13360",-- 4918
x"12d60",-- 4822
x"114c0",-- 4428
x"123b0",-- 4667
x"12230",-- 4643
x"134e0",-- 4942
x"149b0",-- 5275
x"143b0",-- 5179
x"16410",-- 5697
x"169b0",-- 5787
x"16ea0",-- 5866
x"17bf0",-- 6079
x"18270",-- 6183
x"178c0",-- 6028
x"15830",-- 5507
x"11a10",-- 4513
x"0f220",-- 3874
x"0ceb0",-- 3307
x"0a250",-- 2597
x"08030",-- 2051
x"03950",-- 917
x"005c0",-- 92
x"fbb00",-- -1104
x"f7270",-- -2265
x"f30e0",-- -3314
x"ecdf0",-- -4897
x"e8240",-- -6108
x"e49c0",-- -7012
x"e3160",-- -7402
x"e25b0",-- -7589
x"e13e0",-- -7874
x"dfef0",-- -8209
x"df360",-- -8394
x"de6c0",-- -8596
x"e0c80",-- -7992
x"e3040",-- -7420
x"e4be0",-- -6978
x"e9310",-- -5839
x"ec8e0",-- -4978
x"f0f00",-- -3856
x"f4020",-- -3070
x"f6690",-- -2455
x"f8d70",-- -1833
x"fa9d0",-- -1379
x"fd9e0",-- -610
x"01150",-- 277
x"02550",-- 597
x"03810",-- 897
x"03d60",-- 982
x"03990",-- 921
x"04000",-- 1024
x"02b90",-- 697
x"023e0",-- 574
x"001e0",-- 30
x"fe8a0",-- -374
x"fd400",-- -704
x"fb1f0",-- -1249
x"f9150",-- -1771
x"f7020",-- -2302
x"f52e0",-- -2770
x"f41e0",-- -3042
x"f3bd0",-- -3139
x"f3750",-- -3211
x"f3a60",-- -3162
x"f2bb0",-- -3397
x"f3ba0",-- -3142
x"f4780",-- -2952
x"f5e70",-- -2585
x"f8460",-- -1978
x"fa140",-- -1516
x"fc6e0",-- -914
x"feda0",-- -294
x"01620",-- 354
x"03e00",-- 992
x"05fb0",-- 1531
x"079e0",-- 1950
x"09f40",-- 2548
x"0b2b0",-- 2859
x"0d080",-- 3336
x"0e4f0",-- 3663
x"0f040",-- 3844
x"0f6d0",-- 3949
x"0ef70",-- 3831
x"0f5e0",-- 3934
x"0f3d0",-- 3901
x"0ed20",-- 3794
x"0eea0",-- 3818
x"0e9a0",-- 3738
x"0d420",-- 3394
x"0d540",-- 3412
x"0ca00",-- 3232
x"0c130",-- 3091
x"0cc00",-- 3264
x"0d150",-- 3349
x"0dbc0",-- 3516
x"0df00",-- 3568
x"0e7a0",-- 3706
x"0f9c0",-- 3996
x"10db0",-- 4315
x"113a0",-- 4410
x"121e0",-- 4638
x"11dc0",-- 4572
x"122a0",-- 4650
x"12590",-- 4697
x"11100",-- 4368
x"105a0",-- 4186
x"0ed60",-- 3798
x"0e6d0",-- 3693
x"0c750",-- 3189
x"0ad60",-- 2774
x"09490",-- 2377
x"06a90",-- 1705
x"039f0",-- 927
x"00f90",-- 249
x"fe350",-- -459
x"faaa0",-- -1366
x"f7ee0",-- -2066
x"f50e0",-- -2802
x"f32a0",-- -3286
x"f03e0",-- -4034
x"ee780",-- -4488
x"ece30",-- -4893
x"ead90",-- -5415
x"e9de0",-- -5666
x"e9810",-- -5759
x"e8a00",-- -5984
x"e8990",-- -5991
x"e98d0",-- -5747
x"eacb0",-- -5429
x"ec7d0",-- -4995
x"ed900",-- -4720
x"efa20",-- -4190
x"f0a00",-- -3936
x"f2490",-- -3511
x"f4480",-- -3000
x"f5d50",-- -2603
x"f72f0",-- -2257
x"f8eb0",-- -1813
x"fa750",-- -1419
x"fb830",-- -1149
x"fc4b0",-- -949
x"fc960",-- -874
x"fcc50",-- -827
x"fbfd0",-- -1027
x"fc160",-- -1002
x"fbf80",-- -1032
x"fb570",-- -1193
x"faff0",-- -1281
x"faad0",-- -1363
x"fa1e0",-- -1506
x"f9ae0",-- -1618
x"f95c0",-- -1700
x"f9340",-- -1740
x"f9330",-- -1741
x"f97f0",-- -1665
x"fa170",-- -1513
x"f9f40",-- -1548
x"fa430",-- -1469
x"fab70",-- -1353
x"fb3b0",-- -1221
x"fc390",-- -967
x"fd110",-- -751
x"fe4d0",-- -435
x"ff510",-- -175
x"00570",-- 87
x"01740",-- 372
x"01ef0",-- 495
x"02f40",-- 756
x"03b50",-- 949
x"045f0",-- 1119
x"04ed0",-- 1261
x"05970",-- 1431
x"06300",-- 1584
x"06810",-- 1665
x"07220",-- 1826
x"07590",-- 1881
x"07f60",-- 2038
x"087f0",-- 2175
x"08f70",-- 2295
x"09440",-- 2372
x"099a0",-- 2458
x"0a3c0",-- 2620
x"0b130",-- 2835
x"0b530",-- 2899
x"0bd10",-- 3025
x"0c730",-- 3187
x"0c900",-- 3216
x"0d470",-- 3399
x"0d760",-- 3446
x"0de20",-- 3554
x"0df00",-- 3568
x"0e7d0",-- 3709
x"0ed60",-- 3798
x"0ef20",-- 3826
x"0f290",-- 3881
x"0ed60",-- 3798
x"0e820",-- 3714
x"0dc10",-- 3521
x"0d920",-- 3474
x"0d590",-- 3417
x"0d150",-- 3349
x"0cb90",-- 3257
x"0bf10",-- 3057
x"0b0b0",-- 2827
x"09ce0",-- 2510
x"08410",-- 2113
x"06930",-- 1683
x"04a90",-- 1193
x"02e10",-- 737
x"01090",-- 265
x"ff5d0",-- -163
x"fd8f0",-- -625
x"fbd60",-- -1066
x"f9e50",-- -1563
x"f8000",-- -2048
x"f6690",-- -2455
x"f4f00",-- -2832
x"f3c00",-- -3136
x"f2af0",-- -3409
x"f2060",-- -3578
x"f17e0",-- -3714
x"f1250",-- -3803
x"f0cf0",-- -3889
x"f0a30",-- -3933
x"f06b0",-- -3989
x"f0a20",-- -3934
x"f0d00",-- -3888
x"f14f0",-- -3761
x"f1fc0",-- -3588
x"f2930",-- -3437
x"f3560",-- -3242
x"f3720",-- -3214
x"f3830",-- -3197
x"f3520",-- -3246
x"f35c0",-- -3236
x"f3700",-- -3216
x"f3680",-- -3224
x"f3ac0",-- -3156
x"f4050",-- -3067
x"f4480",-- -3000
x"f4cd0",-- -2867
x"f5600",-- -2720
x"f5bd0",-- -2627
x"f6480",-- -2488
x"f6cb0",-- -2357
x"f75b0",-- -2213
x"f8080",-- -2040
x"f8df0",-- -1825
x"f9920",-- -1646
x"fa750",-- -1419
x"fb420",-- -1214
x"fc210",-- -991
x"fd340",-- -716
x"fe350",-- -459
x"ff5d0",-- -163
x"00670",-- 103
x"015b0",-- 347
x"02430",-- 579
x"02f90",-- 761
x"03b30",-- 947
x"046c0",-- 1132
x"050e0",-- 1294
x"05b20",-- 1458
x"063e0",-- 1598
x"06e00",-- 1760
x"07710",-- 1905
x"07e70",-- 2023
x"08550",-- 2133
x"08cc0",-- 2252
x"09360",-- 2358
x"09950",-- 2453
x"09ea0",-- 2538
x"0a3c0",-- 2620
x"0aae0",-- 2734
x"0af90",-- 2809
x"0b330",-- 2867
x"0b680",-- 2920
x"0b7b0",-- 2939
x"0b920",-- 2962
x"0bab0",-- 2987
x"0ba10",-- 2977
x"0bab0",-- 2987
x"0b9f0",-- 2975
x"0b9a0",-- 2970
x"0bb20",-- 2994
x"0bb80",-- 3000
x"0bab0",-- 2987
x"0bcc0",-- 3020
x"0bab0",-- 2987
x"0b860",-- 2950
x"0b710",-- 2929
x"0b380",-- 2872
x"0b330",-- 2867
x"0b2b0",-- 2859
x"0b130",-- 2835
x"0a9b0",-- 2715
x"0a170",-- 2583
x"09900",-- 2448
x"090d0",-- 2317
x"082a0",-- 2090
x"07260",-- 1830
x"05d50",-- 1493
x"04260",-- 1062
x"027d0",-- 637
x"00bb0",-- 187
x"ff360",-- -202
x"fd810",-- -639
x"fc190",-- -999
x"fad90",-- -1319
x"f9b70",-- -1609
x"f89e0",-- -1890
x"f7700",-- -2192
x"f6490",-- -2487
x"f5360",-- -2762
x"f4870",-- -2937
x"f4160",-- -3050
x"f3ef0",-- -3089
x"f3d40",-- -3116
x"f3c70",-- -3129
x"f3950",-- -3179
x"f35b0",-- -3237
x"f3200",-- -3296
x"f2f50",-- -3339
x"f2d50",-- -3371
x"f2cf0",-- -3377
x"f30b0",-- -3317
x"f3470",-- -3257
x"f3970",-- -3177
x"f3c90",-- -3127
x"f3d10",-- -3119
x"f3cf0",-- -3121
x"f3e80",-- -3096
x"f4280",-- -3032
x"f4580",-- -2984
x"f4b20",-- -2894
x"f53e0",-- -2754
x"f5c70",-- -2617
x"f66c0",-- -2452
x"f7340",-- -2252
x"f7df0",-- -2081
x"f8670",-- -1945
x"f91a0",-- -1766
x"fa070",-- -1529
x"fae40",-- -1308
x"fbce0",-- -1074
x"fcc60",-- -826
x"fda40",-- -604
x"fe6e0",-- -402
x"ff5d0",-- -163
x"00340",-- 52
x"00f50",-- 245
x"01900",-- 400
x"022f0",-- 559
x"02cd0",-- 717
x"03650",-- 869
x"040d0",-- 1037
x"04940",-- 1172
x"051d0",-- 1309
x"05990",-- 1433
x"061b0",-- 1563
x"068e0",-- 1678
x"06ef0",-- 1775
x"07240",-- 1828
x"07440",-- 1860
x"074f0",-- 1871
x"074e0",-- 1870
x"07770",-- 1911
x"07770",-- 1911
x"076d0",-- 1901
x"076a0",-- 1898
x"07710",-- 1905
x"076a0",-- 1898
x"07620",-- 1890
x"07510",-- 1873
x"072c0",-- 1836
x"07120",-- 1810
x"07180",-- 1816
x"073b0",-- 1851
x"073b0",-- 1851
x"07440",-- 1860
x"07420",-- 1858
x"07420",-- 1858
x"072b0",-- 1835
x"072b0",-- 1835
x"07150",-- 1813
x"06eb0",-- 1771
x"06d10",-- 1745
x"06a90",-- 1705
x"066c0",-- 1644
x"061c0",-- 1564
x"05d50",-- 1493
x"057c0",-- 1404
x"05490",-- 1353
x"04fc0",-- 1276
x"04cd0",-- 1229
x"04930",-- 1171
x"045d0",-- 1117
x"04260",-- 1062
x"03df0",-- 991
x"039a0",-- 922
x"03350",-- 821
x"02e10",-- 737
x"025f0",-- 607
x"01e00",-- 480
x"01420",-- 322
x"00b60",-- 182
x"001b0",-- 27
x"ff760",-- -138
x"fedc0",-- -292
x"fe3e0",-- -450
x"fdbf0",-- -577
x"fd290",-- -727
x"fcaf0",-- -849
x"fc350",-- -971
x"fbea0",-- -1046
x"fb9a0",-- -1126
x"fb570",-- -1193
x"fb1f0",-- -1249
x"fad20",-- -1326
x"fa930",-- -1389
x"fa410",-- -1471
x"f9fb0",-- -1541
x"f9ae0",-- -1618
x"f9790",-- -1671
x"f92f0",-- -1745
x"f8e40",-- -1820
x"f8a20",-- -1886
x"f8710",-- -1935
x"f8490",-- -1975
x"f8210",-- -2015
x"f7fd0",-- -2051
x"f7db0",-- -2085
x"f7b50",-- -2123
x"f7b00",-- -2128
x"f7c70",-- -2105
x"f7d00",-- -2096
x"f7f30",-- -2061
x"f8230",-- -2013
x"f85c0",-- -1956
x"f89d0",-- -1891
x"f8f20",-- -1806
x"f93e0",-- -1730
x"f9a10",-- -1631
x"fa070",-- -1529
x"fa6e0",-- -1426
x"fada0",-- -1318
x"fb4c0",-- -1204
x"fbd50",-- -1067
x"fc480",-- -952
x"fcdc0",-- -804
x"fd5e0",-- -674
x"fddd0",-- -547
x"fe570",-- -425
x"fede0",-- -290
x"ff510",-- -175
x"ffd60",-- -42
x"00340",-- 52
x"00a30",-- 163
x"01290",-- 297
x"01900",-- 400
x"01fd0",-- 509
x"02520",-- 594
x"02b90",-- 697
x"030e0",-- 782
x"03720",-- 882
x"03bf0",-- 959
x"041b0",-- 1051
x"04690",-- 1129
x"04a50",-- 1189
x"04e80",-- 1256
x"051a0",-- 1306
x"05540",-- 1364
x"057b0",-- 1403
x"05990",-- 1433
x"05b20",-- 1458
x"05bf0",-- 1471
x"05c70",-- 1479
x"05c70",-- 1479
x"05c40",-- 1476
x"05b50",-- 1461
x"05990",-- 1433
x"05830",-- 1411
x"05600",-- 1376
x"05400",-- 1344
x"05120",-- 1298
x"04de0",-- 1246
x"04a50",-- 1189
x"045a0",-- 1114
x"04200",-- 1056
x"03e90",-- 1001
x"03ad0",-- 941
x"03680",-- 872
x"03290",-- 809
x"02d20",-- 722
x"02910",-- 657
x"02610",-- 609
x"02190",-- 537
x"01e50",-- 485
x"01a90",-- 425
x"01720",-- 370
x"01420",-- 322
x"01100",-- 272
x"00e60",-- 230
x"00b60",-- 182
x"00850",-- 133
x"00710",-- 113
x"00440",-- 68
x"001e0",-- 30
x"fffe0",-- -2
x"ffdb0",-- -37
x"ffb50",-- -75
x"ff8f0",-- -113
x"ff790",-- -135
x"ff630",-- -157
x"ff510",-- -175
x"ff310",-- -207
x"ff070",-- -249
x"fedc0",-- -292
x"feb70",-- -329
x"fe9b0",-- -357
x"fe760",-- -394
x"fe500",-- -432
x"fe350",-- -459
x"fe0a0",-- -502
x"fde50",-- -539
x"fdc40",-- -572
x"fd9c0",-- -612
x"fd800",-- -640
x"fd680",-- -664
x"fd4e0",-- -690
x"fd440",-- -700
x"fd1b0",-- -741
x"fd090",-- -759
x"fd070",-- -761
x"fd060",-- -762
x"fd010",-- -767
x"fcf50",-- -779
x"fd010",-- -767
x"fced0",-- -787
x"fce30",-- -797
x"fcee0",-- -786
x"fce40",-- -796
x"fce40",-- -796
x"fced0",-- -787
x"fcf00",-- -784
x"fcfc0",-- -772
x"fd070",-- -761
x"fd240",-- -732
x"fd2f0",-- -721
x"fd3a0",-- -710
x"fd5d0",-- -675
x"fd7b0",-- -645
x"fd9c0",-- -612
x"fdc10",-- -575
x"fdee0",-- -530
x"fe080",-- -504
x"fe410",-- -447
x"fe730",-- -397
x"fea00",-- -352
x"fed20",-- -302
x"fef00",-- -272
x"ff380",-- -200
x"ff670",-- -153
x"ff9f0",-- -97
x"fff10",-- -15
x"00320",-- 50
x"00690",-- 105
x"00a20",-- 162
x"00e40",-- 228
x"01220",-- 290
x"016a0",-- 362
x"019a0",-- 410
x"01cc0",-- 460
x"01f60",-- 502
x"02260",-- 550
x"024d0",-- 589
x"027a0",-- 634
x"02930",-- 659
x"02ac0",-- 684
x"02ca0",-- 714
x"02cc0",-- 716
x"02d90",-- 729
x"02db0",-- 731
x"02e60",-- 742
x"02e80",-- 744
x"02ea0",-- 746
x"02e80",-- 744
x"02d70",-- 727
x"02ca0",-- 714
x"02b10",-- 689
x"02a00",-- 672
x"028f0",-- 655
x"02800",-- 640
x"02550",-- 597
x"02430",-- 579
x"02260",-- 550
x"02050",-- 517
x"01f60",-- 502
x"01c10",-- 449
x"018f0",-- 399
x"01620",-- 354
x"01490",-- 329
x"010d0",-- 269
x"00eb0",-- 235
x"00be0",-- 190
x"007a0",-- 122
x"00580",-- 88
x"00250",-- 37
x"fff80",-- -8
x"ffbc0",-- -68
x"ff8d0",-- -115
x"ff5d0",-- -163
x"ff3a0",-- -198
x"ff0c0",-- -244
x"feed0",-- -275
x"feca0",-- -310
x"feac0",-- -340
x"fe960",-- -362
x"fe800",-- -384
x"fe780",-- -392
x"fe710",-- -399
x"fe5a0",-- -422
x"fe490",-- -439
x"fe440",-- -444
x"fe440",-- -444
x"fe500",-- -432
x"fe530",-- -429
x"fe500",-- -432
x"fe550",-- -427
x"fe5f0",-- -417
x"fe5c0",-- -420
x"fe690",-- -407
x"fe7d0",-- -387
x"fe850",-- -379
x"fe9e0",-- -354
x"fea20",-- -350
x"feb20",-- -334
x"febe0",-- -322
x"fecf0",-- -305
x"feeb0",-- -277
x"fef80",-- -264
x"ff060",-- -250
x"ff100",-- -240
x"ff1f0",-- -225
x"ff260",-- -218
x"ff420",-- -190
x"ff5d0",-- -163
x"ff720",-- -142
x"ff900",-- -112
x"ffad0",-- -83
x"ffd30",-- -45
x"ffd80",-- -40
x"fff10",-- -15
x"fffe0",-- -2
x"00160",-- 22
x"003a0",-- 58
x"00460",-- 70
x"006b0",-- 107
x"006e0",-- 110
x"00800",-- 128
x"00960",-- 150
x"009d0",-- 157
x"00a70",-- 167
x"00af0",-- 175
x"00be0",-- 190
x"00ca0",-- 202
x"00c50",-- 197
x"00c80",-- 200
x"00d90",-- 217
x"00d90",-- 217
x"00e10",-- 225
x"00e40",-- 228
x"00f70",-- 247
x"00f90",-- 249
x"00f70",-- 247
x"00f90",-- 249
x"01030",-- 259
x"01090",-- 265
x"01060",-- 262
x"01150",-- 277
x"010d0",-- 269
x"01100",-- 272
x"01130",-- 275
x"01120",-- 274
x"010b0",-- 267
x"00f90",-- 249
x"00f50",-- 245
x"00eb0",-- 235
x"00eb0",-- 235
x"00dc0",-- 220
x"00d20",-- 210
x"00be0",-- 190
x"00bc0",-- 188
x"00b20",-- 178
x"00a00",-- 160
x"00ac0",-- 172
x"00800",-- 128
x"00730",-- 115
x"00530",-- 83
x"00320",-- 50
x"002b0",-- 43
x"00160",-- 22
x"fffe0",-- -2
x"fff10",-- -15
x"ffdd0",-- -35
x"ffd00",-- -48
x"ffbf0",-- -65
x"ffab0",-- -85
x"ffad0",-- -83
x"ff970",-- -105
x"ff8a0",-- -118
x"ff860",-- -122
x"ff860",-- -122
x"ff8a0",-- -118
x"ff710",-- -143
x"ff620",-- -158
x"ff590",-- -167
x"ff540",-- -172
x"ff490",-- -183
x"ff400",-- -192
x"ff3b0",-- -197
x"ff2b0",-- -213
x"ff1f0",-- -225
x"ff100",-- -240
x"ff070",-- -249
x"fef50",-- -267
x"fef20",-- -270
x"fede0",-- -290
x"fecf0",-- -305
x"fed50",-- -299
x"fed70",-- -297
x"fecf0",-- -305
x"fec60",-- -314
x"febb0",-- -325
x"febe0",-- -322
x"febb0",-- -325
x"fec00",-- -320
x"fed40",-- -300
x"fedc0",-- -292
x"fef50",-- -267
x"fefa0",-- -262
x"ff070",-- -249
x"ff180",-- -232
x"ff110",-- -239
x"ff260",-- -218
x"ff3d0",-- -195
x"ff3b0",-- -197
x"ff450",-- -187
x"ff560",-- -170
x"ff680",-- -152
x"ff7c0",-- -132
x"ff8a0",-- -118
x"ff8d0",-- -115
x"ff9e0",-- -98
x"ffb30",-- -77
x"ffc70",-- -57
x"ffd00",-- -48
x"ffe40",-- -28
x"fffe0",-- -2
x"00110",-- 17
x"002b0",-- 43
x"003a0",-- 58
x"004d0",-- 77
x"005f0",-- 95
x"00710",-- 113
x"00760",-- 118
x"008a0",-- 138
x"009d0",-- 157
x"00b20",-- 178
x"00b40",-- 180
x"00b70",-- 183
x"00c00",-- 192
x"00c30",-- 195
x"00d90",-- 217
x"00e80",-- 232
x"00e40",-- 228
x"00e40",-- 228
x"00ef0",-- 239
x"00f40",-- 244
x"00f00",-- 240
x"00f70",-- 247
x"00fe0",-- 254
x"00eb0",-- 235
x"00e40",-- 228
x"00ed0",-- 237
x"00e80",-- 232
x"00e10",-- 225
x"00cb0",-- 203
x"00bc0",-- 188
x"00b40",-- 180
x"00b20",-- 178
x"00aa0",-- 170
x"00a30",-- 163
x"008a0",-- 138
x"00840",-- 132
x"00780",-- 120
x"005d0",-- 93
x"005c0",-- 92
x"004e0",-- 78
x"00390",-- 57
x"00280",-- 40
x"001e0",-- 30
x"000f0",-- 15
x"fffb0",-- -5
x"fff40",-- -12
x"ffef0",-- -17
x"ffdd0",-- -35
x"ffd50",-- -43
x"ffdf0",-- -33
x"ffc20",-- -62
x"ffae0",-- -82
x"ffb50",-- -75
x"ffb70",-- -73
x"ffb20",-- -78
x"ff940",-- -108
x"ff8f0",-- -113
x"ff830",-- -125
x"ff8b0",-- -117
x"ff800",-- -128
x"ff720",-- -142
x"ff720",-- -142
x"ff650",-- -155
x"ff580",-- -168
x"ff5d0",-- -163
x"ff510",-- -175
x"ff490",-- -183
x"ff4a0",-- -182
x"ff470",-- -185
x"ff510",-- -175
x"ff530",-- -173
x"ff530",-- -173
x"ff590",-- -167
x"ff580",-- -168
x"ff580",-- -168
x"ff6a0",-- -150
x"ff600",-- -160
x"ff740",-- -140
x"ff7e0",-- -130
x"ff7e0",-- -130
x"ff8d0",-- -115
x"ff830",-- -125
x"ff920",-- -110
x"ff950",-- -107
x"ff900",-- -112
x"ff9c0",-- -100
x"ff9e0",-- -98
x"ffa10",-- -95
x"ffa90",-- -87
x"ffb70",-- -73
x"ff9f0",-- -97
x"ffb20",-- -78
x"ffba0",-- -70
x"ffc40",-- -60
x"ffd30",-- -45
x"ffd50",-- -43
x"ffe20",-- -30
x"ffe70",-- -25
x"fff10",-- -15
x"fff60",-- -10
x"fff10",-- -15
x"ffe20",-- -30
x"fff40",-- -12
x"fffb0",-- -5
x"fff30",-- -13
x"00030",-- 3
x"00030",-- 3
x"fffe0",-- -2
x"001e0",-- 30
x"001c0",-- 28
x"00250",-- 37
x"00280",-- 40
x"00170",-- 23
x"00260",-- 38
x"00300",-- 48
x"003e0",-- 62
x"00300",-- 48
x"00440",-- 68
x"003f0",-- 63
x"00320",-- 50
x"00670",-- 103
x"003c0",-- 60
x"00530",-- 83
x"00410",-- 65
x"003a0",-- 58
x"00800",-- 128
x"001e0",-- 30
x"004b0",-- 75
x"005c0",-- 92
x"00370",-- 55
x"004b0",-- 75
x"003c0",-- 60
x"00160",-- 22
x"00440",-- 68
x"003e0",-- 62
x"002f0",-- 47
x"00480",-- 72
x"00200",-- 32
x"004d0",-- 77
x"003f0",-- 63
x"00250",-- 37
x"003a0",-- 58
x"00320",-- 50
x"00370",-- 55
x"00250",-- 37
x"00370",-- 55
x"00260",-- 38
x"000c0",-- 12
x"00170",-- 23
x"00260",-- 38
x"00170",-- 23
x"00000",-- 0
x"00110",-- 17
x"ffe20",-- -30
x"00000",-- 0
x"fffb0",-- -5
x"ffec0",-- -20
x"ffea0",-- -22
x"fff60",-- -10
x"ffdb0",-- -37
x"ffbf0",-- -65
x"ffe20",-- -30
x"ffbd0",-- -67
x"ffce0",-- -50
x"00000",-- 0
x"ffea0",-- -22
x"ffd10",-- -47
x"ffe20",-- -30
x"fff10",-- -15
x"ffa90",-- -87
x"000f0",-- 15
x"ffc20",-- -62
x"ffdf0",-- -33
x"00000",-- 0
x"ffe20",-- -30
x"fffb0",-- -5
x"ffcb0",-- -53
x"00210",-- 33
x"ffe40",-- -28
x"001b0",-- 27
x"ffb80",-- -72
x"00160",-- 22
x"fff80",-- -8
x"ffd80",-- -40
x"001e0",-- 30
x"ffdd0",-- -35
x"000f0",-- 15
x"ffe00",-- -32
x"00080",-- 8
x"00050",-- 5
x"ffdf0",-- -33
x"00110",-- 17
x"00280",-- 40
x"ffe20",-- -30
x"003f0",-- 63
x"fff80",-- -8
x"00160",-- 22
x"00110",-- 17
x"00410",-- 65
x"001e0",-- 30
x"ffdf0",-- -33
x"00410",-- 65
x"00020",-- 2
x"00480",-- 72
x"ffd30",-- -45
x"004e0",-- 78
x"00070",-- 7
x"002b0",-- 43
x"000a0",-- 10
x"00190",-- 25
x"00080",-- 8
x"ffe40",-- -28
x"004d0",-- 77
x"ffc20",-- -62
x"00340",-- 52
x"00070",-- 7
x"00160",-- 22
x"ffe20",-- -30
x"00280",-- 40
x"fff80",-- -8
x"00620",-- 98
x"ffdb0",-- -37
x"ffa80",-- -88
x"00280",-- 40
x"ff630",-- -157
x"fff10",-- -15
x"ffa90",-- -87
x"ffe20",-- -30
x"ff990",-- -103
x"ff9e0",-- -98
x"ffb20",-- -78
x"ff8a0",-- -118
x"ff600",-- -160
x"ff210",-- -223
x"ffa10",-- -95
x"ff6d0",-- -147
x"00570",-- 87
x"ffdd0",-- -35
x"00210",-- 33
x"fff90",-- -7
x"ffdf0",-- -33
x"008f0",-- 143
x"ffa60",-- -90
x"003a0",-- 58
x"00530",-- 83
x"fff10",-- -15
x"003f0",-- 63
x"00430",-- 67
x"00120",-- 18
x"008c0",-- 140
x"ffe20",-- -30
x"000c0",-- 12
x"00520",-- 82
x"ffc40",-- -60
x"004b0",-- 75
x"ff270",-- -217
x"ffba0",-- -70
x"00300",-- 48
x"ff5b0",-- -165
x"00170",-- 23
x"fffb0",-- -5
x"ff710",-- -143
x"fffd0",-- -3
x"ffdf0",-- -33
x"ff4a0",-- -182
x"ffee0",-- -18
x"002b0",-- 43
x"00280",-- 40
x"fed90",-- -295
x"00690",-- 105
x"ff9c0",-- -100
x"00110",-- 17
x"00000",-- 0
x"ffe20",-- -30
x"001e0",-- 30
x"ff510",-- -175
x"00960",-- 150
x"ff620",-- -158
x"fff80",-- -8
x"ffea0",-- -22
x"fffb0",-- -5
x"00070",-- 7
x"fffb0",-- -5
x"000d0",-- 13
x"ff9c0",-- -100
x"008c0",-- 140
x"008f0",-- 143
x"ffdd0",-- -35
x"000d0",-- 13
x"fff40",-- -12
x"001e0",-- 30
x"00110",-- 17
x"00280",-- 40
x"00480",-- 72
x"ff8f0",-- -113
x"00fa0",-- 250
x"005a0",-- 90
x"ffe00",-- -32
x"00530",-- 83
x"00440",-- 68
x"00000",-- 0
x"ffdb0",-- -37
x"00a80",-- 168
x"000f0",-- 15
x"009d0",-- 157
x"ff5e0",-- -162
x"001e0",-- 30
x"00250",-- 37
x"008f0",-- 143
x"00210",-- 33
x"ff6d0",-- -147
x"00e30",-- 227
x"ffa60",-- -90
x"00d20",-- 210
x"ffb70",-- -73
x"00000",-- 0
x"fffb0",-- -5
x"00200",-- 32
x"ffa60",-- -90
x"00940",-- 148
x"00110",-- 17
x"ffe00",-- -32
x"00210",-- 33
x"fffd0",-- -3
x"007d0",-- 125
x"ffce0",-- -50
x"00e80",-- 232
x"ff210",-- -223
x"00850",-- 133
x"ffad0",-- -83
x"00cb0",-- 203
x"ff5e0",-- -162
x"00140",-- 20
x"00000",-- 0
x"ff990",-- -103
x"01620",-- 354
x"fe7a0",-- -390
x"01210",-- 289
x"ffbf0",-- -65
x"00670",-- 103
x"ff9c0",-- -100
x"00210",-- 33
x"ffab0",-- -85
x"ffce0",-- -50
x"00460",-- 70
x"ff2c0",-- -212
x"00a30",-- 163
x"fef70",-- -265
x"008c0",-- 140
x"ff6a0",-- -150
x"00530",-- 83
x"ff4f0",-- -177
x"ffce0",-- -50
x"ffae0",-- -82
x"00280",-- 40
x"fff80",-- -8
x"feca0",-- -310
x"00700",-- 112
x"ffc20",-- -62
x"ffe50",-- -27
x"00350",-- 53
x"ffdd0",-- -35
x"ffe00",-- -32
x"fff10",-- -15
x"ffe50",-- -27
x"00550",-- 85
x"ff530",-- -173
x"ffdb0",-- -37
x"ff7c0",-- -132
x"004e0",-- 78
x"ff790",-- -135
x"00370",-- 55
x"000c0",-- 12
x"ff940",-- -108
x"002d0",-- 45
x"ffe50",-- -27
x"00940",-- 148
x"ff8f0",-- -113
x"ff620",-- -158
x"00780",-- 120
x"ff240",-- -220
x"00c00",-- 192
x"ff9f0",-- -97
x"00500",-- 80
x"ff6d0",-- -147
x"ffea0",-- -22
x"00570",-- 87
x"ff270",-- -217
x"007b0",-- 123
x"ffc60",-- -58
x"ff3d0",-- -195
x"01060",-- 262
x"fe710",-- -399
x"00e80",-- 232
x"00750",-- 117
x"fef30",-- -269
x"015b0",-- 347
x"ff590",-- -167
x"00170",-- 23
x"ff600",-- -160
x"00000",-- 0
x"000f0",-- 15
x"ffa30",-- -93
x"00460",-- 70
x"00200",-- 32
x"00660",-- 102
x"ffd60",-- -42
x"00160",-- 22
x"ff9a0",-- -102
x"00000",-- 0
x"ff940",-- -108
x"ffc20",-- -62
x"00440",-- 68
x"ff860",-- -122
x"00250",-- 37
x"00530",-- 83
x"00660",-- 102
x"004b0",-- 75
x"003a0",-- 58
x"ffb80",-- -72
x"ffce0",-- -50
x"ff5d0",-- -163
x"00f70",-- 247
x"ff830",-- -125
x"00cb0",-- 203
x"ff680",-- -152
x"00230",-- 35
x"00700",-- 112
x"ff580",-- -168
x"010b0",-- 267
x"fe980",-- -360
x"01880",-- 392
x"fecf0",-- -305
x"00140",-- 20
x"00b10",-- 177
x"fea80",-- -344
x"00a70",-- 167
x"ffc70",-- -57
x"000f0",-- 15
x"ff6a0",-- -150
x"01540",-- 340
x"ff450",-- -187
x"00d90",-- 217
x"fedf0",-- -289
x"00780",-- 120
x"ff720",-- -142
x"ff010",-- -255
x"01150",-- 277
x"fe700",-- -400
x"00d70",-- 215
x"ff400",-- -192
x"010d0",-- 269
x"ff010",-- -255
x"00c00",-- 192
x"ff530",-- -173
x"008c0",-- 140
x"ffec0",-- -20
x"fec10",-- -319
x"00ff0",-- 255
x"ff0e0",-- -242
x"00980",-- 152
x"ff2b0",-- -213
x"ffd60",-- -42
x"ffa60",-- -90
x"00af0",-- 175
x"ff490",-- -183
x"00a00",-- 160
x"fff10",-- -15
x"fea00",-- -352
x"005a0",-- 90
x"009e0",-- 158
x"009d0",-- 157
x"ff510",-- -175
x"00eb0",-- 235
x"ff2b0",-- -213
x"fffb0",-- -5
x"002f0",-- 47
x"002f0",-- 47
x"003a0",-- 58
x"00370",-- 55
x"00050",-- 5
x"00230",-- 35
x"00af0",-- 175
x"ffa30",-- -93
x"ffdf0",-- -33
x"00a00",-- 160
x"ff3b0",-- -197
x"00a00",-- 160
x"ff8a0",-- -118
x"01350",-- 309
x"005a0",-- 90
x"ff180",-- -232
x"01a30",-- 419
x"fe390",-- -455
x"01bd0",-- 445
x"ff9f0",-- -97
x"ffa90",-- -87
x"01040",-- 260
x"fe990",-- -359
x"00d40",-- 212
x"ff4e0",-- -178
x"00e60",-- 230
x"ffc90",-- -55
x"00750",-- 117
x"00300",-- 48
x"00230",-- 35
x"ffc60",-- -58
x"ff580",-- -168
x"01950",-- 405
x"ff670",-- -153
x"005f0",-- 95
x"ff600",-- -160
x"00760",-- 118
x"00320",-- 50
x"ff8a0",-- -118
x"00080",-- 8
x"00940",-- 148
x"ff6a0",-- -150
x"ffb80",-- -72
x"00e40",-- 228
x"ffc60",-- -58
x"00e40",-- 228
x"002b0",-- 43
x"ff790",-- -135
x"00a50",-- 165
x"ffba0",-- -70
x"00d00",-- 208
x"ffbd0",-- -67
x"ff630",-- -157
x"00a70",-- 167
x"febe0",-- -322
x"00c00",-- 192
x"006b0",-- 107
x"ffda0",-- -38
x"010d0",-- 269
x"ff440",-- -188
x"ffbf0",-- -65
x"00410",-- 65
x"ffec0",-- -20
x"ff3a0",-- -198
x"01360",-- 310
x"feb60",-- -330
x"012e0",-- 302
x"ff920",-- -110
x"003e0",-- 62
x"00250",-- 37
x"febe0",-- -322
x"01ce0",-- 462
x"feca0",-- -310
x"ffbf0",-- -65
x"00550",-- 85
x"ff310",-- -207
x"00800",-- 128
x"00a30",-- 163
x"ff510",-- -175
x"00890",-- 137
x"ff530",-- -173
x"ffce0",-- -50
x"ffea0",-- -22
x"002b0",-- 43
x"00080",-- 8
x"ff2e0",-- -210
x"00280",-- 40
x"fff30",-- -13
x"00c80",-- 200
x"ffb30",-- -77
x"ffe20",-- -30
x"00aa0",-- 170
x"fdf60",-- -522
x"011a0",-- 282
x"ffa30",-- -93
x"ff290",-- -215
x"00f50",-- 245
x"fec50",-- -315
x"001c0",-- 28
x"ffad0",-- -83
x"008f0",-- 143
x"01580",-- 344
x"fd8d0",-- -627
x"01e70",-- 487
x"ff350",-- -203
x"fe980",-- -360
x"02120",-- 530
x"fe210",-- -479
x"01090",-- 265
x"00480",-- 72
x"ff6f0",-- -145
x"00190",-- 25
x"fff90",-- -7
x"000c0",-- 12
x"01540",-- 340
x"ff540",-- -172
x"ff5d0",-- -163
x"003e0",-- 62
x"fff80",-- -8
x"ff8a0",-- -118
x"ff110",-- -239
x"00320",-- 50
x"ff070",-- -249
x"014e0",-- 334
x"ff290",-- -215
x"01710",-- 369
x"fe850",-- -379
x"00a80",-- 168
x"006c0",-- 108
x"fe8e0",-- -370
x"01f40",-- 500
x"fd940",-- -620
x"01c90",-- 457
x"fead0",-- -339
x"ffc90",-- -55
x"01100",-- 272
x"ff180",-- -232
x"00d50",-- 213
x"ffa30",-- -93
x"002f0",-- 47
x"00eb0",-- 235
x"fff80",-- -8
x"ff240",-- -220
x"011c0",-- 284
x"fef70",-- -265
x"00260",-- 38
x"00b10",-- 177
x"feb10",-- -335
x"02320",-- 562
x"fe170",-- -489
x"01f90",-- 505
x"fe980",-- -360
x"00690",-- 105
x"012c0",-- 300
x"fe9e0",-- -354
x"00c80",-- 200
x"feda0",-- -294
x"00050",-- 5
x"ff770",-- -137
x"00430",-- 67
x"ffc90",-- -55
x"ffd50",-- -43
x"00d00",-- 208
x"ff6c0",-- -148
x"01150",-- 277
x"fee10",-- -287
x"ff3b0",-- -197
x"01a60",-- 422
x"fda40",-- -604
x"01180",-- 280
x"004b0",-- 75
x"fdc70",-- -569
x"02960",-- 662
x"ff5d0",-- -163
x"00870",-- 135
x"013d0",-- 317
x"fe080",-- -504
x"01b50",-- 437
x"ff110",-- -239
x"ff0e0",-- -242
x"01ce0",-- 462
x"fe1b0",-- -485
x"00af0",-- 175
x"00410",-- 65
x"ffa30",-- -93
x"00490",-- 73
x"fee30",-- -285
x"008c0",-- 140
x"006b0",-- 107
x"fff10",-- -15
x"000f0",-- 15
x"fff60",-- -10
x"ffad0",-- -83
x"ffe90",-- -23
x"fe620",-- -414
x"ff950",-- -107
x"02520",-- 594
x"fee10",-- -287
x"00700",-- 112
x"00000",-- 0
x"ff4a0",-- -182
x"009e0",-- 158
x"ffd80",-- -40
x"ff900",-- -112
x"00960",-- 150
x"fd2e0",-- -722
x"02020",-- 514
x"00e40",-- 228
x"fdce0",-- -562
x"02350",-- 565
x"fea00",-- -352
x"01090",-- 265
x"febb0",-- -325
x"ffe50",-- -27
x"007f0",-- 127
x"ff3b0",-- -197
x"ffba0",-- -70
x"00cb0",-- 203
x"004e0",-- 78
x"ff290",-- -215
x"00080",-- 8
x"007d0",-- 125
x"feeb0",-- -277
x"00610",-- 97
x"00460",-- 70
x"000d0",-- 13
x"ffd00",-- -48
x"ffbf0",-- -65
x"02200",-- 544
x"fd440",-- -700
x"02390",-- 569
x"fdcb0",-- -565
x"01a60",-- 422
x"fe9e0",-- -354
x"ff8a0",-- -118
x"01b00",-- 432
x"fe2a0",-- -470
x"024d0",-- 589
x"fd3d0",-- -707
x"02ed0",-- 749
x"fdee0",-- -530
x"00280",-- 40
x"00890",-- 137
x"fda90",-- -599
x"027f0",-- 639
x"fe000",-- -512
x"01420",-- 322
x"fe2d0",-- -467
x"00d20",-- 210
x"ff630",-- -157
x"01620",-- 354
x"fe0a0",-- -502
x"011a0",-- 282
x"fefd0",-- -259
x"fefa0",-- -262
x"00bc0",-- 188
x"fe3a0",-- -454
x"03ae0",-- 942
x"fbd80",-- -1064
x"03920",-- 914
x"fcf70",-- -777
x"03420",-- 834
x"fc890",-- -887
x"01350",-- 309
x"00610",-- 97
x"fe1b0",-- -485
x"04f50",-- 1269
x"f98b0",-- -1653
x"06c20",-- 1730
x"f9f90",-- -1543
x"01df0",-- 479
x"01a90",-- 425
x"fe280",-- -472
x"02120",-- 530
x"fb3d0",-- -1219
x"03fd0",-- 1021
x"fe250",-- -475
x"01450",-- 325
x"fe870",-- -377
x"01900",-- 400
x"fe0f0",-- -497
x"ffa60",-- -90
x"01b00",-- 432
x"fd160",-- -746
x"00eb0",-- 235
x"ff0b0",-- -245
x"01620",-- 354
x"ff270",-- -217
x"00b70",-- 183
x"fee40",-- -284
x"ff210",-- -223
x"02170",-- 535
x"fe570",-- -425
x"028a0",-- 650
x"fd110",-- -751
x"01420",-- 322
x"007a0",-- 122
x"ff950",-- -107
x"016c0",-- 364
x"fed70",-- -297
x"00ac0",-- 172
x"fd240",-- -732
x"02cd0",-- 717
x"fe6b0",-- -405
x"00170",-- 23
x"00fc0",-- 252
x"fe8a0",-- -374
x"026e0",-- 622
x"fd1d0",-- -739
x"02570",-- 599
x"fe3a0",-- -454
x"00c50",-- 197
x"001b0",-- 27
x"fdec0",-- -532
x"02170",-- 535
x"fe300",-- -464
x"006b0",-- 107
x"01ba0",-- 442
x"00670",-- 103
x"ffec0",-- -20
x"004e0",-- 78
x"fd360",-- -714
x"01ea0",-- 490
x"fd8f0",-- -625
x"035d0",-- 861
x"fd130",-- -749
x"01970",-- 407
x"ff7c0",-- -132
x"ff4c0",-- -180
x"033d0",-- 829
x"fdae0",-- -594
x"01ce0",-- 462
x"fe0f0",-- -497
x"ff3b0",-- -197
x"00250",-- 37
x"00f00",-- 240
x"02140",-- 532
x"fecd0",-- -307
x"015e0",-- 350
x"fcd70",-- -809
x"01f80",-- 504
x"00230",-- 35
x"fe410",-- -447
x"03310",-- 817
x"fb880",-- -1144
x"022b0",-- 555
x"fd8b0",-- -629
x"02f40",-- 756
x"fc3c0",-- -964
x"00d50",-- 213
x"01e90",-- 489
x"fc5c0",-- -932
x"04520",-- 1106
x"fc500",-- -944
x"03770",-- 887
x"fddb0",-- -549
x"01310",-- 305
x"00d50",-- 213
x"fe940",-- -364
x"ffc20",-- -62
x"01620",-- 354
x"00e30",-- 227
x"ff620",-- -158
x"02c10",-- 705
x"fe990",-- -359
x"ffc70",-- -57
x"010d0",-- 269
x"ff580",-- -168
x"ffc60",-- -58
x"01150",-- 277
x"fd6c0",-- -660
x"01800",-- 384
x"fdb20",-- -590
x"00c30",-- 195
x"fde00",-- -544
x"fcb20",-- -846
x"04820",-- 1154
x"fcb40",-- -844
x"01770",-- 375
x"01260",-- 294
x"fe080",-- -504
x"02e00",-- 736
x"fe9d0",-- -355
x"fff10",-- -15
x"ffa10",-- -95
x"fea00",-- -352
x"02fe0",-- 766
x"fee40",-- -284
x"ff010",-- -255
x"02f70",-- 759
x"00890",-- 137
x"00780",-- 120
x"ff490",-- -183
x"011d0",-- 285
x"ffd00",-- -48
x"fe850",-- -379
x"ffc40",-- -60
x"fed00",-- -304
x"00170",-- 23
x"003e0",-- 62
x"ffb20",-- -78
x"00990",-- 153
x"00250",-- 37
x"00490",-- 73
x"00a50",-- 165
x"fe230",-- -477
x"01f40",-- 500
x"fea50",-- -347
x"fcd00",-- -816
x"00550",-- 85
x"00700",-- 112
x"fbc70",-- -1081
x"02520",-- 594
x"00c50",-- 197
x"fff10",-- -15
x"fdb50",-- -587
x"012e0",-- 302
x"01cb0",-- 459
x"fc710",-- -911
x"01f40",-- 500
x"fed70",-- -297
x"000a0",-- 10
x"00460",-- 70
x"02030",-- 515
x"fde70",-- -537
x"02250",-- 549
x"fff10",-- -15
x"ff710",-- -143
x"01540",-- 340
x"000c0",-- 12
x"01290",-- 297
x"fd990",-- -615
x"00530",-- 83
x"00d40",-- 212
x"ffa90",-- -87
x"ff070",-- -249
x"031a0",-- 794
x"fd0e0",-- -754
x"01990",-- 409
x"fee90",-- -279
x"ff350",-- -203
x"01a80",-- 424
x"fd2a0",-- -726
x"02ca0",-- 714
x"fb7c0",-- -1156
x"02120",-- 530
x"fe070",-- -505
x"00210",-- 33
x"ffd30",-- -45
x"feac0",-- -340
x"01580",-- 344
x"fe730",-- -397
x"03220",-- 802
x"fd720",-- -654
x"00800",-- 128
x"fea20",-- -350
x"03c10",-- 961
x"fcd90",-- -807
x"03420",-- 834
x"014f0",-- 335
x"fdfe0",-- -514
x"02be0",-- 702
x"fbef0",-- -1041
x"02de0",-- 734
x"fce40",-- -796
x"04440",-- 1092
x"fe570",-- -425
x"01620",-- 354
x"01b30",-- 435
x"fa700",-- -1424
x"05810",-- 1409
x"fa9e0",-- -1378
x"03b20",-- 946
x"01420",-- 322
x"fd3a0",-- -710
x"02550",-- 597
x"fc870",-- -889
x"00160",-- 22
x"ff110",-- -239
x"01740",-- 372
x"ffc20",-- -62
x"fe700",-- -400
x"02110",-- 529
x"fe170",-- -489
x"01970",-- 407
x"fce40",-- -796
x"00ff0",-- 255
x"00370",-- 55
x"fef20",-- -270
x"04030",-- 1027
x"ff860",-- -122
x"fe6b0",-- -405
x"00e40",-- 228
x"ff2b0",-- -213
x"023c0",-- 572
x"ff6d0",-- -147
x"fd7b0",-- -645
x"05310",-- 1329
x"fbf60",-- -1034
x"04f90",-- 1273
x"fde00",-- -544
x"00460",-- 70
x"000a0",-- 10
x"fc2d0",-- -979
x"02350",-- 565
x"fe570",-- -425
x"013b0",-- 315
x"fe8c0",-- -372
x"040d0",-- 1037
x"fd2a0",-- -726
x"fe660",-- -410
x"00d70",-- 215
x"ff9c0",-- -100
x"013d0",-- 317
x"fecf0",-- -305
x"04710",-- 1137
x"fc8e0",-- -882
x"02c30",-- 707
x"fe760",-- -394
x"fff90",-- -7
x"00df0",-- 223
x"fc160",-- -1002
x"038a0",-- 906
x"fdfb0",-- -517
x"ffb20",-- -78
x"017b0",-- 379
x"fd8d0",-- -627
x"ff1f0",-- -225
x"00990",-- 153
x"02f20",-- 754
x"ff4f0",-- -177
x"ff3f0",-- -193
x"03400",-- 832
x"fc390",-- -967
x"03130",-- 787
x"fd310",-- -719
x"01510",-- 337
x"fee90",-- -279
x"00500",-- 80
x"02120",-- 530
x"fc200",-- -992
x"06780",-- 1656
x"f7e70",-- -2073
x"04c50",-- 1221
x"fea80",-- -344
x"000f0",-- 15
x"03300",-- 816
x"012b0",-- 299
x"ff010",-- -255
x"ffe50",-- -27
x"020a0",-- 522
x"f9c60",-- -1594
x"03880",-- 904
x"fc230",-- -989
x"04f40",-- 1268
x"ff310",-- -207
x"00280",-- 40
x"01a60",-- 422
x"fc3c0",-- -964
x"05770",-- 1399
x"fae30",-- -1309
x"ffc20",-- -62
x"ff760",-- -138
x"00fe0",-- 254
x"fd990",-- -615
x"036c0",-- 876
x"fe0d0",-- -499
x"fd180",-- -744
x"046c0",-- 1132
x"fa940",-- -1388
x"06c20",-- 1730
x"f9a30",-- -1629
x"05940",-- 1428
x"fbee0",-- -1042
x"00f50",-- 245
x"001e0",-- 30
x"fc030",-- -1021
x"050e0",-- 1294
x"fcdf0",-- -801
x"00250",-- 37
x"01400",-- 320
x"030e0",-- 782
x"f9610",-- -1695
x"06500",-- 1616
x"f8d20",-- -1838
x"02260",-- 550
x"fd1a0",-- -742
x"01380",-- 312
x"01a90",-- 425
x"f9540",-- -1708
x"0c5f0",-- 3167
x"f3b50",-- -3147
x"07100",-- 1808
x"ff330",-- -205
x"ff420",-- -190
x"ffe50",-- -27
x"fe570",-- -425
x"06a40",-- 1700
x"f5950",-- -2667
x"07ad0",-- 1965
x"01e40",-- 484
x"f94c0",-- -1716
x"013f0",-- 319
x"025c0",-- 604
x"ff710",-- -143
x"00160",-- 22
x"004e0",-- 78
x"038b0",-- 907
x"fc990",-- -871
x"002f0",-- 47
x"ff490",-- -183
x"fcc30",-- -829
x"02670",-- 615
x"002d0",-- 45
x"05c70",-- 1479
x"fcf20",-- -782
x"fc5c0",-- -932
x"07920",-- 1938
x"f8cd0",-- -1843
x"00bb0",-- 187
x"06710",-- 1649
x"f95b0",-- -1701
x"04fc0",-- 1276
x"f9420",-- -1726
x"04760",-- 1142
x"fdfe0",-- -514
x"fa710",-- -1423
x"05ad0",-- 1453
x"fe370",-- -457
x"fdb30",-- -589
x"00dc0",-- 220
x"02f70",-- 759
x"f7d50",-- -2091
x"04750",-- 1141
x"fbf10",-- -1039
x"ffa80",-- -88
x"ff790",-- -135
x"fe890",-- -375
x"03300",-- 816
x"fe020",-- -510
x"03560",-- 854
x"fb940",-- -1132
x"fd090",-- -759
x"04ae0",-- 1198
x"fbc20",-- -1086
x"ff220",-- -222
x"07770",-- 1911
x"fa440",-- -1468
x"04c70",-- 1223
x"fe000",-- -512
x"fcd00",-- -816
x"009d0",-- 157
x"ff5d0",-- -163
x"01760",-- 374
x"fe120",-- -494
x"066b0",-- 1643
x"faaa0",-- -1366
x"03ba0",-- 954
x"ff950",-- -107
x"fe250",-- -475
x"014f0",-- 335
x"00dc0",-- 220
x"01510",-- 337
x"00000",-- 0
x"fdf30",-- -525
x"024e0",-- 590
x"fbc60",-- -1082
x"ffa10",-- -95
x"02390",-- 569
x"f9fe0",-- -1538
x"07350",-- 1845
x"ffea0",-- -22
x"01030",-- 259
x"ffc90",-- -55
x"fe570",-- -425
x"febe0",-- -322
x"fd240",-- -732
x"023c0",-- 572
x"01620",-- 354
x"fe700",-- -400
x"01220",-- 290
x"fd740",-- -652
x"02070",-- 519
x"ff770",-- -137
x"fce10",-- -799
x"07220",-- 1826
x"fbd30",-- -1069
x"063c0",-- 1596
x"ff580",-- -168
x"fddb0",-- -549
x"04690",-- 1129
x"fcd90",-- -807
x"066c0",-- 1644
x"fe780",-- -392
x"033b0",-- 827
x"01170",-- 279
x"fcc50",-- -827
x"04820",-- 1154
x"fb920",-- -1134
x"03240",-- 804
x"fa3c0",-- -1476
x"02390",-- 569
x"03010",-- 769
x"fa350",-- -1483
x"07ef0",-- 2031
x"f8110",-- -2031
x"026c0",-- 620
x"fd4f0",-- -689
x"01620",-- 354
x"ffc90",-- -55
x"fc3f0",-- -961
x"04dc0",-- 1244
x"f59f0",-- -2657
x"08210",-- 2081
x"fadc0",-- -1316
x"fe850",-- -379
x"01a60",-- 422
x"fa2a0",-- -1494
x"03810",-- 897
x"fd850",-- -635
x"fe3e0",-- -450
x"01f90",-- 505
x"fd680",-- -664
x"007a0",-- 122
x"05060",-- 1286
x"f9f10",-- -1551
x"06710",-- 1649
x"fbe90",-- -1047
x"ffdb0",-- -37
x"05580",-- 1368
x"fce60",-- -794
x"03740",-- 884
x"ffbd0",-- -67
x"00e80",-- 232
x"00700",-- 112
x"03bd0",-- 957
x"fffd0",-- -3
x"00980",-- 152
x"006c0",-- 108
x"01fb0",-- 507
x"02870",-- 647
x"fc6e0",-- -914
x"04f20",-- 1266
x"fed40",-- -300
x"fe340",-- -460
x"059f0",-- 1439
x"fde20",-- -542
x"03a80",-- 936
x"fdd10",-- -559
x"ffd50",-- -43
x"04340",-- 1076
x"fad70",-- -1321
x"00410",-- 65
x"01ec0",-- 492
x"fa120",-- -1518
x"00870",-- 135
x"01290",-- 297
x"fe910",-- -367
x"017c0",-- 380
x"fd5b0",-- -677
x"00190",-- 25
x"fd8b0",-- -629
x"ffab0",-- -85
x"00260",-- 38
x"fce30",-- -797
x"019c0",-- 412
x"fe070",-- -505
x"01c90",-- 457
x"fd6f0",-- -657
x"00960",-- 150
x"fe990",-- -359
x"01ae0",-- 430
x"ff800",-- -128
x"fe890",-- -375
x"04ae0",-- 1198
x"fb2f0",-- -1233
x"019f0",-- 415
x"fd770",-- -649
x"ffa60",-- -90
x"fff40",-- -12
x"ff3a0",-- -198
x"01970",-- 407
x"fd220",-- -734
x"039f0",-- 927
x"fd2e0",-- -722
x"fd8d0",-- -627
x"ff170",-- -233
x"fdbd0",-- -579
x"00d40",-- 212
x"00e10",-- 225
x"00fe0",-- 254
x"00990",-- 153
x"fd530",-- -685
x"fc890",-- -887
x"04660",-- 1126
x"fdd10",-- -559
x"000f0",-- 15
x"01b00",-- 432
x"fe780",-- -392
x"013f0",-- 319
x"ffb80",-- -72
x"fe580",-- -424
x"feaa0",-- -342
x"01bf0",-- 447
x"fe8e0",-- -370
x"04e10",-- 1249
x"ff860",-- -122
x"00170",-- 23
x"ffea0",-- -22
x"fae30",-- -1309
x"034c0",-- 844
x"fecb0",-- -309
x"037c0",-- 892
x"fe4e0",-- -434
x"ffdf0",-- -33
x"04260",-- 1062
x"fc0a0",-- -1014
x"02460",-- 582
x"fe340",-- -460
x"fdbc0",-- -580
x"04f50",-- 1269
x"00850",-- 133
x"02160",-- 534
x"015d0",-- 349
x"fd2c0",-- -724
x"fdab0",-- -597
x"01310",-- 305
x"01970",-- 407
x"02670",-- 615
x"00980",-- 152
x"ff790",-- -135
x"02a70",-- 679
x"fe760",-- -394
x"ffdd0",-- -35
x"00e30",-- 227
x"fde00",-- -544
x"02f00",-- 752
x"01450",-- 325
x"01210",-- 289
x"00500",-- 80
x"fc980",-- -872
x"ff770",-- -137
x"ff950",-- -107
x"00e10",-- 225
x"00cd0",-- 205
x"00210",-- 33
x"005c0",-- 92
x"ffce0",-- -50
x"fe460",-- -442
x"ff800",-- -128
x"fe7f0",-- -385
x"ff670",-- -153
x"01a90",-- 425
x"01740",-- 372
x"001b0",-- 27
x"fe730",-- -397
x"fee80",-- -280
x"fe610",-- -415
x"ff860",-- -122
x"00480",-- 72
x"022f0",-- 559
x"00780",-- 120
x"ff040",-- -252
x"ff4e0",-- -178
x"fee60",-- -282
x"ff990",-- -103
x"ff1c0",-- -228
x"03210",-- 801
x"00570",-- 87
x"02120",-- 530
x"01e50",-- 485
x"fc2d0",-- -979
x"01100",-- 272
x"ff8a0",-- -118
x"ff860",-- -122
x"000f0",-- 15
x"01170",-- 279
x"00530",-- 83
x"fecd0",-- -307
x"ffbf0",-- -65
x"fe4e0",-- -434
x"ffe70",-- -25
x"ff5d0",-- -163
x"ffdf0",-- -33
x"01a10",-- 417
x"00800",-- 128
x"fd360",-- -714
x"fd3b0",-- -709
x"fff10",-- -15
x"fe570",-- -425
x"00410",-- 65
x"00320",-- 50
x"00a30",-- 163
x"01d30",-- 467
x"fff40",-- -12
x"ffec0",-- -20
x"002f0",-- 47
x"ff680",-- -152
x"00ef0",-- 239
x"02db0",-- 731
x"007f0",-- 127
x"02b90",-- 697
x"ff680",-- -152
x"00340",-- 52
x"ff8d0",-- -115
x"017c0",-- 380
x"03090",-- 777
x"00280",-- 40
x"029e0",-- 670
x"010e0",-- 270
x"00280",-- 40
x"fed40",-- -300
x"ff8b0",-- -117
x"ff150",-- -235
x"ffcc0",-- -52
x"01770",-- 375
x"01490",-- 329
x"000c0",-- 12
x"fd510",-- -687
x"fdc90",-- -567
x"fef70",-- -265
x"fff10",-- -15
x"00af0",-- 175
x"fea20",-- -350
x"000c0",-- 12
x"ff210",-- -223
x"fe930",-- -365
x"fffb0",-- -5
x"fd160",-- -746
x"007a0",-- 122
x"008a0",-- 138
x"015b0",-- 347
x"02550",-- 597
x"fef50",-- -267
x"fe850",-- -379
x"ff940",-- -108
x"002a0",-- 42
x"01e90",-- 489
x"02490",-- 585
x"fd8b0",-- -629
x"ff530",-- -173
x"fe5f0",-- -417
x"ff680",-- -152
x"010d0",-- 269
x"fed70",-- -297
x"ff510",-- -175
x"fee60",-- -282
x"ffbc0",-- -68
x"005a0",-- 90
x"fe960",-- -362
x"fccb0",-- -821
x"fe690",-- -407
x"00480",-- 72
x"01f80",-- 504
x"02030",-- 515
x"00170",-- 23
x"fecf0",-- -305
x"ffab0",-- -85
x"01ec0",-- 492
x"03010",-- 769
x"032e0",-- 814
x"02990",-- 665
x"01420",-- 322
x"024b0",-- 587
x"02640",-- 612
x"01580",-- 344
x"01d30",-- 467
x"00df0",-- 223
x"007a0",-- 122
x"02500",-- 592
x"01470",-- 327
x"ff070",-- -249
x"fdb50",-- -587
x"fde70",-- -537
x"ff330",-- -205
x"008a0",-- 138
x"00570",-- 87
x"fd990",-- -615
x"fcc60",-- -826
x"fcfc0",-- -772
x"fdd10",-- -559
x"fe820",-- -382
x"fe300",-- -464
x"fd470",-- -697
x"fec80",-- -312
x"feb90",-- -327
x"fed40",-- -300
x"fe320",-- -462
x"fd630",-- -669
x"feda0",-- -294
x"00030",-- 3
x"01260",-- 294
x"00e60",-- 230
x"ffa30",-- -93
x"feb70",-- -329
x"ffbd0",-- -67
x"01770",-- 375
x"023f0",-- 575
x"01900",-- 400
x"01540",-- 340
x"01220",-- 290
x"01040",-- 260
x"01680",-- 360
x"014f0",-- 335
x"00de0",-- 222
x"013f0",-- 319
x"02300",-- 560
x"029d0",-- 669
x"01e00",-- 480
x"019a0",-- 410
x"007a0",-- 122
x"00e40",-- 228
x"01940",-- 404
x"025a0",-- 602
x"00cb0",-- 203
x"00800",-- 128
x"ffe00",-- -32
x"ff2e0",-- -210
x"00110",-- 17
x"ff400",-- -192
x"ffae0",-- -82
x"ff590",-- -167
x"ff150",-- -235
x"ff3d0",-- -195
x"fee90",-- -279
x"fe070",-- -505
x"fdfb0",-- -517
x"fe260",-- -474
x"fdd50",-- -555
x"fea80",-- -344
x"fe000",-- -512
x"fcf70",-- -777
x"fd9f0",-- -609
x"fe030",-- -509
x"fec50",-- -315
x"fea70",-- -345
x"feda0",-- -294
x"fe780",-- -392
x"fed40",-- -300
x"ff5b0",-- -165
x"ffc60",-- -58
x"fff60",-- -10
x"000c0",-- 12
x"006c0",-- 108
x"00f90",-- 249
x"01860",-- 390
x"01710",-- 369
x"023e0",-- 574
x"02190",-- 537
x"01d00",-- 464
x"017c0",-- 380
x"02660",-- 614
x"02b70",-- 695
x"02e30",-- 739
x"03120",-- 786
x"02120",-- 530
x"021c0",-- 540
x"019c0",-- 412
x"01e40",-- 484
x"01920",-- 402
x"00f20",-- 242
x"00c00",-- 192
x"ffdf0",-- -33
x"ff920",-- -110
x"ff3b0",-- -197
x"fe700",-- -400
x"fe140",-- -492
x"fd600",-- -672
x"fd470",-- -697
x"fd3d0",-- -707
x"fcfc0",-- -772
x"fcf20",-- -782
x"fd1a0",-- -742
x"fcfc0",-- -772
x"fd420",-- -702
x"fd600",-- -672
x"fd1d0",-- -739
x"fde90",-- -535
x"fe190",-- -487
x"febe0",-- -322
x"fee80",-- -280
x"ff1f0",-- -225
x"ff070",-- -249
x"ff470",-- -185
x"00690",-- 105
x"00760",-- 118
x"01650",-- 357
x"012c0",-- 300
x"01880",-- 392
x"01620",-- 354
x"019e0",-- 414
x"01790",-- 377
x"01f10",-- 497
x"01fd0",-- 509
x"01cb0",-- 459
x"01fd0",-- 509
x"01360",-- 310
x"01560",-- 342
x"00bc0",-- 188
x"01180",-- 280
x"00cb0",-- 203
x"00cf0",-- 207
x"00670",-- 103
x"00160",-- 22
x"ff9e0",-- -98
x"ff260",-- -218
x"ff560",-- -170
x"fee10",-- -287
x"ff400",-- -192
x"febe0",-- -322
x"fea70",-- -345
x"fe980",-- -360
x"fe120",-- -494
x"fe4d0",-- -435
x"fe140",-- -492
x"fe410",-- -447
x"fe940",-- -364
x"fed70",-- -297
x"fea50",-- -347
x"feda0",-- -294
x"fe8f0",-- -369
x"ff1c0",-- -228
x"ff560",-- -170
x"ffdb0",-- -37
x"fff10",-- -15
x"00320",-- 50
x"00700",-- 112
x"001b0",-- 27
x"00a30",-- 163
x"00c60",-- 198
x"01180",-- 280
x"01350",-- 309
x"017c0",-- 380
x"01860",-- 390
x"017b0",-- 379
x"01770",-- 375
x"018f0",-- 399
x"01740",-- 372
x"019a0",-- 410
x"01900",-- 400
x"012c0",-- 300
x"010e0",-- 270
x"00cb0",-- 203
x"008f0",-- 143
x"00750",-- 117
x"00430",-- 67
x"00230",-- 35
x"ffc70",-- -57
x"ffb00",-- -80
x"ff7b0",-- -133
x"ff240",-- -220
x"ff010",-- -255
x"fefa0",-- -262
x"feda0",-- -294
x"fea50",-- -347
x"feb40",-- -332
x"fe800",-- -384
x"fe9e0",-- -354
x"feaa0",-- -342
x"feb20",-- -334
x"febc0",-- -324
x"fed00",-- -304
x"fef30",-- -269
x"ff1c0",-- -228
x"ff400",-- -192
x"ff810",-- -127
x"ffa40",-- -92
x"ffba0",-- -70
x"ffdb0",-- -37
x"00000",-- 0
x"00200",-- 32
x"004b0",-- 75
x"00b90",-- 185
x"00a00",-- 160
x"00d50",-- 213
x"009b0",-- 155
x"00bc0",-- 188
x"009d0",-- 157
x"00eb0",-- 235
x"00ef0",-- 239
x"00c50",-- 197
x"01030",-- 259
x"00990",-- 153
x"00af0",-- 175
x"00760",-- 118
x"007b0",-- 123
x"00480",-- 72
x"00610",-- 97
x"00410",-- 65
x"00200",-- 32
x"fffb0",-- -5
x"ffb80",-- -72
x"ffbc0",-- -68
x"ff8a0",-- -118
x"ffc10",-- -63
x"ff900",-- -112
x"ff740",-- -140
x"ff5d0",-- -163
x"ff4e0",-- -178
x"ff4a0",-- -182
x"ff530",-- -173
x"ff5e0",-- -162
x"ff530",-- -173
x"ff4e0",-- -178
x"ff560",-- -170
x"ff710",-- -143
x"ff5d0",-- -163
x"ff8a0",-- -118
x"ff4f0",-- -177
x"ffb20",-- -78
x"ffb50",-- -75
x"ffd50",-- -43
x"00260",-- 38
x"fff40",-- -12
x"003e0",-- 62
x"000c0",-- 12
x"00610",-- 97
x"00520",-- 82
x"00620",-- 98
x"00580",-- 88
x"00700",-- 112
x"00730",-- 115
x"00620",-- 98
x"006b0",-- 107
x"00280",-- 40
x"005f0",-- 95
x"005d0",-- 93
x"00730",-- 115
x"005c0",-- 92
x"002b0",-- 43
x"00250",-- 37
x"fffb0",-- -5
x"002b0",-- 43
x"00000",-- 0
x"002b0",-- 43
x"ffea0",-- -22
x"ffe40",-- -28
x"ffe40",-- -28
x"ffae0",-- -82
x"ffc40",-- -60
x"ff9a0",-- -102
x"ffe70",-- -25
x"ffa90",-- -87
x"ffd10",-- -47
x"ffb00",-- -80
x"ff940",-- -108
x"ffb00",-- -80
x"ff8a0",-- -118
x"fff30",-- -13
x"ffd50",-- -43
x"ffec0",-- -20
x"ffe20",-- -30
x"ffd60",-- -42
x"ffec0",-- -20
x"ffdb0",-- -37
x"ffea0",-- -22
x"fff60",-- -10
x"00080",-- 8
x"00120",-- 18
x"00000",-- 0
x"fff80",-- -8
x"fffe0",-- -2
x"00030",-- 3
x"00120",-- 18
x"00110",-- 17
x"002f0",-- 47
x"00020",-- 2
x"002d0",-- 45
x"00000",-- 0
x"00050",-- 5
x"00250",-- 37
x"000c0",-- 12
x"00120",-- 18
x"fffe0",-- -2
x"00110",-- 17
x"fff80",-- -8
x"00110",-- 17
x"ffe50",-- -27
x"ffee0",-- -18
x"ffe70",-- -25
x"fff90",-- -7
x"fff30",-- -13
x"ffc60",-- -58
x"fff40",-- -12
x"ffa60",-- -90
x"ffd50",-- -43
x"ffc20",-- -62
x"ffbf0",-- -65
x"ffc90",-- -55
x"ffbd0",-- -67
x"ffc70",-- -57
x"ffb20",-- -78
x"ffd80",-- -40
x"ffc90",-- -55
x"ffb80",-- -72
x"ffe50",-- -27
x"ffd80",-- -40
x"ffee0",-- -18
x"fff10",-- -15
x"ffe00",-- -32
x"ffda0",-- -38
x"00030",-- 3
x"00020",-- 2
x"00050",-- 5
x"00070",-- 7
x"000c0",-- 12
x"000f0",-- 15
x"00140",-- 20
x"000f0",-- 15
x"00070",-- 7
x"001b0",-- 27
x"001c0",-- 28
x"00340",-- 52
x"00200",-- 32
x"00120",-- 18
x"00020",-- 2
x"000a0",-- 10
x"fffe0",-- -2
x"00050",-- 5
x"00000",-- 0
x"fffd0",-- -3
x"fff10",-- -15
x"ffe70",-- -25
x"ffdf0",-- -33
x"ffc90",-- -55
x"ffd80",-- -40
x"ffc60",-- -58
x"ffea0",-- -22
x"ffd80",-- -40
x"ffb50",-- -75
x"ffe20",-- -30
x"ffc20",-- -62
x"ffda0",-- -38
x"ffbf0",-- -65
x"ffd30",-- -45
x"ffdd0",-- -35
x"ffbc0",-- -68
x"ffe70",-- -25
x"ffc90",-- -55
x"ffe20",-- -30
x"ffd30",-- -45
x"ffe20",-- -30
x"ffe50",-- -27
x"ffd10",-- -47
x"fff60",-- -10
x"ffce0",-- -50
x"00070",-- 7
x"ffe90",-- -23
x"ffe40",-- -28
x"fff90",-- -7
x"ffda0",-- -38
x"00000",-- 0
x"ffe50",-- -27
x"00000",-- 0
x"ffee0",-- -18
x"ffdb0",-- -37
x"ffe90",-- -23
x"ffe90",-- -23
x"ffd10",-- -47
x"ffd60",-- -42
x"ffdf0",-- -33
x"ffd10",-- -47
x"ffe20",-- -30
x"ffd50",-- -43
x"ffdf0",-- -33
x"ffc20",-- -62
x"ffdd0",-- -35
x"ffd80",-- -40
x"ffe00",-- -32
x"ffe20",-- -30
x"ffdb0",-- -37
x"ffdd0",-- -35
x"ffda0",-- -38
x"ffdd0",-- -35
x"ffea0",-- -22
x"ffea0",-- -22
x"ffee0",-- -18
x"ffdd0",-- -35
x"fff40",-- -12
x"ffef0",-- -17
x"ffe90",-- -23
x"fff40",-- -12
x"ffce0",-- -50
x"00000",-- 0
x"ffda0",-- -38
x"fff60",-- -10
x"fff10",-- -15
x"ffee0",-- -18
x"00050",-- 5
x"ffe40",-- -28
x"00120",-- 18
x"fffb0",-- -5
x"000c0",-- 12
x"00070",-- 7
x"00030",-- 3
x"002b0",-- 43
x"00000",-- 0
x"001e0",-- 30
x"00000",-- 0
x"00160",-- 22
x"00200",-- 32
x"00200",-- 32
x"00260",-- 38
x"00000",-- 0
x"00370",-- 55
x"000f0",-- 15
x"00300",-- 48
x"00320",-- 50
x"00170",-- 23
x"003a0",-- 58
x"00210",-- 33
x"00320",-- 50
x"00280",-- 40
x"00280",-- 40
x"00300",-- 48
x"001e0",-- 30
x"002f0",-- 47
x"00280",-- 40
x"00230",-- 35
x"00320",-- 50
x"001c0",-- 28
x"00280",-- 40
x"001c0",-- 28
x"00390",-- 57
x"00340",-- 52
x"00350",-- 53
x"00490",-- 73
x"00350",-- 53
x"00500",-- 80
x"003a0",-- 58
x"002b0",-- 43
x"00370",-- 55
x"00370",-- 55
x"00390",-- 57
x"002a0",-- 42
x"00430",-- 67
x"002f0",-- 47
x"00250",-- 37
x"002d0",-- 45
x"00280",-- 40
x"002a0",-- 42
x"00370",-- 55
x"00300",-- 48
x"001c0",-- 28
x"00200",-- 32
x"00200",-- 32
x"00210",-- 33
x"001b0",-- 27
x"000f0",-- 15
x"00190",-- 25
x"000a0",-- 10
x"001b0",-- 27
x"00120",-- 18
x"00120",-- 18
x"00030",-- 3
x"000f0",-- 15
x"001b0",-- 27
x"fff90",-- -7
x"001b0",-- 27
x"000a0",-- 10
x"00050",-- 5
x"fff40",-- -12
x"000d0",-- 13
x"00030",-- 3
x"00000",-- 0
x"001c0",-- 28
x"fff80",-- -8
x"001b0",-- 27
x"00020",-- 2
x"00080",-- 8
x"fffd0",-- -3
x"00020",-- 2
x"000a0",-- 10
x"fffd0",-- -3
x"00210",-- 33
x"fff10",-- -15
x"00160",-- 22
x"00080",-- 8
x"00070",-- 7
x"00050",-- 5
x"00030",-- 3
x"00050",-- 5
x"fffb0",-- -5
x"00160",-- 22
x"00120",-- 18
x"00020",-- 2
x"00000",-- 0
x"00080",-- 8
x"00020",-- 2
x"00020",-- 2
x"fff30",-- -13
x"fffb0",-- -5
x"ffef0",-- -17
x"00000",-- 0
x"00030",-- 3
x"fff30",-- -13
x"00030",-- 3
x"ffea0",-- -22
x"ffe70",-- -25
x"fff80",-- -8
x"fff10",-- -15
x"ffea0",-- -22
x"fff10",-- -15
x"ffef0",-- -17
x"ffe90",-- -23
x"fff80",-- -8
x"fff80",-- -8
x"fff30",-- -13
x"fff90",-- -7
x"fff30",-- -13
x"00080",-- 8
x"fff80",-- -8
x"00050",-- 5
x"ffee0",-- -18
x"fffb0",-- -5
x"ffe20",-- -30
x"00000",-- 0
x"fffd0",-- -3
x"ffe20",-- -30
x"fff10",-- -15
x"ffdd0",-- -35
x"00000",-- 0
x"ffe20",-- -30
x"fff40",-- -12
x"ffd30",-- -45
x"ffef0",-- -17
x"fff10",-- -15
x"ffe20",-- -30
x"ffee0",-- -18
x"ffdd0",-- -35
x"fff30",-- -13
x"ffe40",-- -28
x"fff30",-- -13
x"ffdf0",-- -33
x"ffdf0",-- -33
x"ffdf0",-- -33
x"ffd30",-- -45
x"ffdd0",-- -35
x"ffc60",-- -58
x"ffd50",-- -43
x"ffcb0",-- -53
x"ffd80",-- -40
x"ffd00",-- -48
x"ffc90",-- -55
x"ffd80",-- -40
x"ffbf0",-- -65
x"ffdb0",-- -37
x"ffe70",-- -25
x"ffd00",-- -48
x"ffdf0",-- -33
x"ffce0",-- -50
x"ffda0",-- -38
x"ffd10",-- -47
x"ffd60",-- -42
x"ffdb0",-- -37
x"ffd80",-- -40
x"ffea0",-- -22
x"ffcc0",-- -52
x"fff80",-- -8
x"ffdf0",-- -33
x"fff10",-- -15
x"ffe50",-- -27
x"ffd80",-- -40
x"ffea0",-- -22
x"ffc90",-- -55
x"fffb0",-- -5
x"ffdb0",-- -37
x"ffe50",-- -27
x"ffef0",-- -17
x"fff60",-- -10
x"fff40",-- -12
x"ffe70",-- -25
x"fff10",-- -15
x"ffdf0",-- -33
x"fff80",-- -8
x"00000",-- 0
x"00000",-- 0
x"fff30",-- -13
x"fffd0",-- -3
x"fffb0",-- -5
x"fff40",-- -12
x"fff90",-- -7
x"ffe70",-- -25
x"00000",-- 0
x"fffd0",-- -3
x"fff80",-- -8
x"fffb0",-- -5
x"fffb0",-- -5
x"ffef0",-- -17
x"fff80",-- -8
x"00000",-- 0
x"fffb0",-- -5
x"fffe0",-- -2
x"fff90",-- -7
x"fff80",-- -8
x"fff80",-- -8
x"fff80",-- -8
x"fffb0",-- -5
x"00020",-- 2
x"fff40",-- -12
x"00000",-- 0
x"00000",-- 0
x"fffb0",-- -5
x"00030",-- 3
x"ffef0",-- -17
x"fff60",-- -10
x"ffef0",-- -17
x"fffd0",-- -3
x"fff10",-- -15
x"ffef0",-- -17
x"fff60",-- -10
x"fff10",-- -15
x"ffee0",-- -18
x"ffef0",-- -17
x"00020",-- 2
x"ffea0",-- -22
x"ffec0",-- -20
x"fff30",-- -13
x"fff80",-- -8
x"fff30",-- -13
x"fff40",-- -12
x"ffee0",-- -18
x"fff10",-- -15
x"00000",-- 0
x"fff90",-- -7
x"fff80",-- -8
x"fff60",-- -10
x"ffe20",-- -30
x"ffee0",-- -18
x"fff80",-- -8
x"ffea0",-- -22
x"ffef0",-- -17
x"ffe50",-- -27
x"fffb0",-- -5
x"ffee0",-- -18
x"ffe50",-- -27
x"fff80",-- -8
x"ffe00",-- -32
x"ffd80",-- -40
x"ffe50",-- -27
x"ffe20",-- -30
x"ffdd0",-- -35
x"ffe20",-- -30
x"ffe20",-- -30
x"ffda0",-- -38
x"ffdb0",-- -37
x"ffef0",-- -17
x"ffdb0",-- -37
x"ffe90",-- -23
x"ffdf0",-- -33
x"ffd30",-- -45
x"ffe40",-- -28
x"ffdf0",-- -33
x"ffce0",-- -50
x"ffd10",-- -47
x"ffce0",-- -50
x"ffd30",-- -45
x"ffd10",-- -47
x"ffd10",-- -47
x"ffd10",-- -47
x"ffc70",-- -57
x"ffce0",-- -50
x"ffc20",-- -62
x"ffdb0",-- -37
x"ffc60",-- -58
x"ffd50",-- -43
x"ffc70",-- -57
x"ffd10",-- -47
x"ffea0",-- -22
x"ffd50",-- -43
x"ffe20",-- -30
x"ffcb0",-- -53
x"ffec0",-- -20
x"ffdb0",-- -37
x"ffe70",-- -25
x"fffd0",-- -3
x"ffea0",-- -22
x"ffe90",-- -23
x"ffdb0",-- -37
x"ffe50",-- -27
x"ffe70",-- -25
x"ffe70",-- -25
x"ffdd0",-- -35
x"ffea0",-- -22
x"ffe20",-- -30
x"ffd60",-- -42
x"ffec0",-- -20
x"ffe20",-- -30
x"ffe40",-- -28
x"ffee0",-- -18
x"ffee0",-- -18
x"fff10",-- -15
x"ffe50",-- -27
x"ffe40",-- -28
x"ffe90",-- -23
x"fff90",-- -7
x"fffe0",-- -2
x"ffec0",-- -20
x"00000",-- 0
x"fff40",-- -12
x"fff40",-- -12
x"ffee0",-- -18
x"fff40",-- -12
x"ffef0",-- -17
x"ffdb0",-- -37
x"fff80",-- -8
x"ffe50",-- -27
x"ffe90",-- -23
x"fff80",-- -8
x"fff40",-- -12
x"ffe50",-- -27
x"ffec0",-- -20
x"ffee0",-- -18
x"ffea0",-- -22
x"fff10",-- -15
x"ffe50",-- -27
x"ffe50",-- -27
x"ffef0",-- -17
x"fff90",-- -7
x"fff30",-- -13
x"ffea0",-- -22
x"fff80",-- -8
x"fff40",-- -12
x"fff10",-- -15
x"ffec0",-- -20
x"fff30",-- -13
x"ffea0",-- -22
x"fff40",-- -12
x"fffb0",-- -5
x"fffe0",-- -2
x"fff10",-- -15
x"00000",-- 0
x"fffe0",-- -2
x"00000",-- 0
x"00140",-- 20
x"00030",-- 3
x"000c0",-- 12
x"00000",-- 0
x"00080",-- 8
x"00000",-- 0
x"00070",-- 7
x"000d0",-- 13
x"00110",-- 17
x"000c0",-- 12
x"00140",-- 20
x"00140",-- 20
x"00020",-- 2
x"00160",-- 22
x"00050",-- 5
x"000f0",-- 15
x"00000",-- 0
x"000c0",-- 12
x"00050",-- 5
x"00020",-- 2
x"00020",-- 2
x"fff90",-- -7
x"000f0",-- 15
x"00020",-- 2
x"00160",-- 22
x"000a0",-- 10
x"000d0",-- 13
x"00070",-- 7
x"00070",-- 7
x"00140",-- 20
x"000a0",-- 10
x"001b0",-- 27
x"00110",-- 17
x"00120",-- 18
x"00170",-- 23
x"00160",-- 22
x"00170",-- 23
x"00170",-- 23
x"00140",-- 20
x"000d0",-- 13
x"00020",-- 2
x"00160",-- 22
x"00160",-- 22
x"000f0",-- 15
x"00140",-- 20
x"00120",-- 18
x"00170",-- 23
x"00120",-- 18
x"001e0",-- 30
x"00160",-- 22
x"001b0",-- 27
x"00160",-- 22
x"000c0",-- 12
x"00160",-- 22
x"000d0",-- 13
x"00080",-- 8
x"00030",-- 3
x"00050",-- 5
x"000c0",-- 12
x"00000",-- 0
x"00050",-- 5
x"00020",-- 2
x"00110",-- 17
x"00020",-- 2
x"00070",-- 7
x"00080",-- 8
x"00000",-- 0
x"00000",-- 0
x"fff30",-- -13
x"00050",-- 5
x"fff40",-- -12
x"00000",-- 0
x"fff40",-- -12
x"00000",-- 0
x"00050",-- 5
x"fff80",-- -8
x"fffd0",-- -3
x"fff40",-- -12
x"00000",-- 0
x"fff10",-- -15
x"00030",-- 3
x"fffe0",-- -2
x"00000",-- 0
x"00070",-- 7
x"fff60",-- -10
x"fff80",-- -8
x"fff80",-- -8
x"00020",-- 2
x"00050",-- 5
x"00050",-- 5
x"00020",-- 2
x"fffb0",-- -5
x"00000",-- 0
x"ffee0",-- -18
x"ffef0",-- -17
x"00000",-- 0
x"00000",-- 0
x"fffb0",-- -5
x"fff80",-- -8
x"00000",-- 0
x"00000",-- 0
x"fff60",-- -10
x"ffee0",-- -18
x"fffb0",-- -5
x"fff80",-- -8
x"ffe90",-- -23
x"fff80",-- -8
x"ffe70",-- -25
x"fff10",-- -15
x"ffe00",-- -32
x"ffea0",-- -22
x"00000",-- 0
x"ffea0",-- -22
x"fff30",-- -13
x"fff10",-- -15
x"fff10",-- -15
x"ffd80",-- -40
x"ffec0",-- -20
x"ffd60",-- -42
x"ffd60",-- -42
x"ffea0",-- -22
x"ffdf0",-- -33
x"ffdb0",-- -37
x"ffd60",-- -42
x"ffdb0",-- -37
x"ffd00",-- -48
x"ffdb0",-- -37
x"ffd30",-- -45
x"ffd50",-- -43
x"ffe00",-- -32
x"ffce0",-- -50
x"ffd80",-- -40
x"ffd00",-- -48
x"ffd10",-- -47
x"ffc70",-- -57
x"ffdb0",-- -37
x"ffd80",-- -40
x"ffd50",-- -43
x"ffdd0",-- -35
x"ffcc0",-- -52
x"ffd80",-- -40
x"ffd80",-- -40
x"ffe50",-- -27
x"ffdd0",-- -35
x"ffe50",-- -27
x"ffe50",-- -27
x"ffee0",-- -18
x"ffea0",-- -22
x"fff10",-- -15
x"ffee0",-- -18
x"ffee0",-- -18
x"00000",-- 0
x"fffb0",-- -5
x"00000",-- 0
x"fffd0",-- -3
x"fffe0",-- -2
x"fff40",-- -12
x"00000",-- 0
x"fff60",-- -10
x"00000",-- 0
x"fff90",-- -7
x"ffea0",-- -22
x"fffe0",-- -2
x"fff40",-- -12
x"fffb0",-- -5
x"fffb0",-- -5
x"00000",-- 0
x"fff40",-- -12
x"00000",-- 0
x"fff90",-- -7
x"fffb0",-- -5
x"00000",-- 0
x"fff40",-- -12
x"00050",-- 5
x"00070",-- 7
x"00070",-- 7
x"00120",-- 18
x"000c0",-- 12
x"00110",-- 17
x"000c0",-- 12
x"00000",-- 0
x"00070",-- 7
x"00000",-- 0
x"00050",-- 5
x"00160",-- 22
x"000d0",-- 13
x"00000",-- 0
x"00000",-- 0
x"000f0",-- 15
x"00070",-- 7
x"00080",-- 8
x"000a0",-- 10
x"000a0",-- 10
x"00050",-- 5
x"000d0",-- 13
x"00080",-- 8
x"00160",-- 22
x"00080",-- 8
x"00080",-- 8
x"00160",-- 22
x"00190",-- 25
x"00080",-- 8
x"000f0",-- 15
x"00170",-- 23
x"000f0",-- 15
x"00120",-- 18
x"00190",-- 25
x"00200",-- 32
x"001c0",-- 28
x"00230",-- 35
x"00140",-- 20
x"00250",-- 37
x"000c0",-- 12
x"00190",-- 25
x"00230",-- 35
x"001c0",-- 28
x"00170",-- 23
x"000d0",-- 13
x"00140",-- 20
x"00080",-- 8
x"00260",-- 38
x"00110",-- 17
x"00110",-- 17
x"001b0",-- 27
x"00160",-- 22
x"00280",-- 40
x"00140",-- 20
x"00160",-- 22
x"00140",-- 20
x"00260",-- 38
x"001b0",-- 27
x"00160",-- 22
x"00160",-- 22
x"00030",-- 3
x"00190",-- 25
x"000a0",-- 10
x"00050",-- 5
x"00070",-- 7
x"00110",-- 17
x"00190",-- 25
x"00120",-- 18
x"00170",-- 23
x"00000",-- 0
x"00020",-- 2
x"00070",-- 7
x"00050",-- 5
x"000c0",-- 12
x"000c0",-- 12
x"00020",-- 2
x"00050",-- 5
x"000c0",-- 12
x"000a0",-- 10
x"00020",-- 2
x"00080",-- 8
x"00000",-- 0
x"fffe0",-- -2
x"00000",-- 0
x"fff40",-- -12
x"fff10",-- -15
x"ffef0",-- -17
x"fffe0",-- -2
x"fff10",-- -15
x"fff60",-- -10
x"ffef0",-- -17
x"ffec0",-- -20
x"fff10",-- -15
x"fff30",-- -13
x"00000",-- 0
x"ffea0",-- -22
x"fff80",-- -8
x"fff90",-- -7
x"fffd0",-- -3
x"fff10",-- -15
x"fffb0",-- -5
x"fff80",-- -8
x"fff60",-- -10
x"fffb0",-- -5
x"fffd0",-- -3
x"00000",-- 0
x"fffe0",-- -2
x"00050",-- 5
x"fffb0",-- -5
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fff30",-- -13
x"00000",-- 0
x"fffe0",-- -2
x"fff90",-- -7
x"fff80",-- -8
x"fff10",-- -15
x"ffec0",-- -20
x"fff30",-- -13
x"00020",-- 2
x"ffee0",-- -18
x"fff90",-- -7
x"fff10",-- -15
x"ffee0",-- -18
x"fff30",-- -13
x"fff60",-- -10
x"ffe50",-- -27
x"ffe00",-- -32
x"ffe50",-- -27
x"ffe50",-- -27
x"ffea0",-- -22
x"ffdb0",-- -37
x"ffea0",-- -22
x"ffd60",-- -42
x"ffd80",-- -40
x"ffda0",-- -38
x"ffdf0",-- -33
x"ffe20",-- -30
x"ffe50",-- -27
x"ffe90",-- -23
x"ffdb0",-- -37
x"ffe20",-- -30
x"ffd50",-- -43
x"ffd80",-- -40
x"ffd80",-- -40
x"ffd60",-- -42
x"ffd50",-- -43
x"ffdb0",-- -37
x"ffd50",-- -43
x"ffda0",-- -38
x"ffe50",-- -27
x"ffdb0",-- -37
x"ffdd0",-- -35
x"ffdd0",-- -35
x"ffce0",-- -50
x"ffd50",-- -43
x"ffe20",-- -30
x"ffcb0",-- -53
x"ffd50",-- -43
x"ffce0",-- -50
x"ffd30",-- -45
x"ffbd0",-- -67
x"ffc90",-- -55
x"ff990",-- -103
x"ffad0",-- -83
x"ff530",-- -173
x"ff540",-- -172
x"fee40",-- -284
x"febe0",-- -322
x"fdea0",-- -534
x"fdbc0",-- -580
x"fb330",-- -1229
x"f5d00",-- -2608
x"fb040",-- -1276
x"00b90",-- 185
x"fe370",-- -457
x"fa6b0",-- -1429
x"f67b0",-- -2437
x"f7790",-- -2183
x"fe570",-- -425
x"00de0",-- 222
x"fe500",-- -432
x"f9b80",-- -1608
x"f8d50",-- -1835
x"ffd10",-- -47
x"06020",-- 1538
x"067d0",-- 1661
x"02930",-- 659
x"00cd0",-- 205
x"06cc0",-- 1740
x"0db20",-- 3506
x"0f540",-- 3924
x"0ca70",-- 3239
x"0b1f0",-- 2847
x"0d1d0",-- 3357
x"0fa40",-- 4004
x"0f650",-- 3941
x"0d9f0",-- 3487
x"0ab60",-- 2742
x"08cc0",-- 2252
x"09060",-- 2310
x"06e50",-- 1765
x"03530",-- 851
x"02480",-- 584
x"023c0",-- 572
x"ff770",-- -137
x"fbc10",-- -1087
x"fada0",-- -1318
x"fad70",-- -1321
x"fa670",-- -1433
x"fa9d0",-- -1379
x"f86e0",-- -1938
x"f5070",-- -2809
x"f6550",-- -2475
x"f98b0",-- -1653
x"f9990",-- -1639
x"f82a0",-- -2006
x"f70e0",-- -2290
x"f6fa0",-- -2310
x"f91d0",-- -1763
x"fc260",-- -986
x"fc2f0",-- -977
x"f9f10",-- -1551
x"f9e20",-- -1566
x"fb790",-- -1159
x"fcf00",-- -784
x"fe140",-- -492
x"fe120",-- -494
x"fd0c0",-- -756
x"fcfc0",-- -772
x"fe660",-- -410
x"ff790",-- -135
x"000a0",-- 10
x"005f0",-- 95
x"00390",-- 57
x"00080",-- 8
x"00910",-- 145
x"01db0",-- 475
x"02f40",-- 756
x"03100",-- 784
x"026b0",-- 619
x"021c0",-- 540
x"025c0",-- 604
x"03670",-- 871
x"04610",-- 1121
x"03ab0",-- 939
x"02610",-- 609
x"01f10",-- 497
x"02580",-- 600
x"02ca0",-- 714
x"03260",-- 806
x"02260",-- 550
x"005d0",-- 93
x"004e0",-- 78
x"00cd0",-- 205
x"00af0",-- 175
x"00520",-- 82
x"ff9f0",-- -97
x"fe7a0",-- -390
x"fdef0",-- -529
x"fea80",-- -344
x"fec80",-- -312
x"fe170",-- -489
x"fe000",-- -512
x"fda40",-- -604
x"fcfc0",-- -772
x"fd9c0",-- -612
x"fe8a0",-- -374
x"fe340",-- -460
x"fe0a0",-- -502
x"fe230",-- -477
x"fde70",-- -537
x"fe760",-- -394
x"ffb80",-- -72
x"ffdf0",-- -33
x"ff440",-- -188
x"ff670",-- -153
x"ffd30",-- -45
x"004b0",-- 75
x"01060",-- 262
x"016a0",-- 362
x"00be0",-- 190
x"00710",-- 113
x"01100",-- 272
x"01740",-- 372
x"01a80",-- 424
x"01990",-- 409
x"013f0",-- 319
x"00c80",-- 200
x"00eb0",-- 235
x"016a0",-- 362
x"01670",-- 359
x"00ff0",-- 255
x"00ad0",-- 173
x"00350",-- 53
x"00050",-- 5
x"00020",-- 2
x"003e0",-- 62
x"ffc60",-- -58
x"ff1a0",-- -230
x"ff350",-- -203
x"fec10",-- -319
x"fefa0",-- -262
x"ff400",-- -192
x"ff0c0",-- -244
x"fea20",-- -350
x"fe850",-- -379
x"fecb0",-- -309
x"feeb0",-- -277
x"fef80",-- -264
x"ff4c0",-- -180
x"fed70",-- -297
x"fea80",-- -344
x"ff040",-- -252
x"ff7e0",-- -130
x"ff310",-- -207
x"fff30",-- -13
x"fde40",-- -540
x"fb620",-- -1182
x"fe340",-- -460
x"009d0",-- 157
x"ff600",-- -160
x"fbcc0",-- -1076
x"f9bc0",-- -1604
x"fb390",-- -1223
x"fe530",-- -429
x"fe1b0",-- -485
x"facd0",-- -1331
x"f7630",-- -2205
x"f8530",-- -1965
x"fbc10",-- -1087
x"fcfc0",-- -772
x"fae40",-- -1308
x"f8a80",-- -1880
x"f98a0",-- -1654
x"fc620",-- -926
x"fe620",-- -414
x"ff8f0",-- -113
x"fff40",-- -12
x"005a0",-- 90
x"03560",-- 854
x"068e0",-- 1678
x"06f70",-- 1783
x"09170",-- 2327
x"0bd50",-- 3029
x"0c2a0",-- 3114
x"0b2e0",-- 2862
x"0c500",-- 3152
x"0eea0",-- 3818
x"12500",-- 4688
x"142c0",-- 5164
x"10c80",-- 4296
x"0c5e0",-- 3166
x"0d950",-- 3477
x"11ee0",-- 4590
x"11e70",-- 4583
x"0cde0",-- 3294
x"07180",-- 1816
x"04700",-- 1136
x"05170",-- 1303
x"06530",-- 1619
x"03e90",-- 1001
x"fe020",-- -510
x"f9130",-- -1773
x"f8610",-- -1951
x"f9df0",-- -1569
x"f9970",-- -1641
x"f77a0",-- -2182
x"f5720",-- -2702
x"f3720",-- -3214
x"f2cf0",-- -3377
x"f5470",-- -2745
x"f7470",-- -2233
x"f6500",-- -2480
x"f5310",-- -2767
x"f5090",-- -2807
x"f51f0",-- -2785
x"f6c30",-- -2365
x"fa640",-- -1436
x"fb1d0",-- -1251
x"f8ad0",-- -1875
x"f8460",-- -1978
x"fa210",-- -1503
x"fc2a0",-- -982
x"fe7f0",-- -385
x"ff270",-- -217
x"fd090",-- -759
x"fbd10",-- -1071
x"fe480",-- -440
x"01630",-- 355
x"02230",-- 547
x"01710",-- 369
x"008f0",-- 143
x"00320",-- 50
x"01c40",-- 452
x"04390",-- 1081
x"05240",-- 1316
x"03720",-- 882
x"02410",-- 577
x"02f70",-- 759
x"03e40",-- 996
x"04d10",-- 1233
x"052c0",-- 1324
x"04200",-- 1056
x"01f80",-- 504
x"01bf0",-- 447
x"03260",-- 806
x"035b0",-- 859
x"026b0",-- 619
x"018f0",-- 399
x"fffe0",-- -2
x"feb40",-- -332
x"fff40",-- -12
x"01080",-- 264
x"ffab0",-- -85
x"fd3d0",-- -707
x"fc440",-- -956
x"fc8f0",-- -881
x"fbb20",-- -1102
x"fc660",-- -922
x"fc390",-- -967
x"fa140",-- -1516
x"f8800",-- -1920
x"f8930",-- -1901
x"f9b50",-- -1611
x"f9ce0",-- -1586
x"f8f80",-- -1800
x"f75e0",-- -2210
x"f6120",-- -2542
x"f6e90",-- -2327
x"f8930",-- -1901
x"f8f70",-- -1801
x"f8500",-- -1968
x"f7570",-- -2217
x"f8250",-- -2011
x"fa120",-- -1518
x"fbad0",-- -1107
x"fce40",-- -796
x"fdae0",-- -594
x"fef00",-- -272
x"00f40",-- 244
x"04a50",-- 1189
x"07b30",-- 1971
x"089d0",-- 2205
x"07300",-- 1840
x"0c630",-- 3171
x"12b10",-- 4785
x"10590",-- 4185
x"0d080",-- 3336
x"0f810",-- 3969
x"13b20",-- 5042
x"158f0",-- 5519
x"18200",-- 6176
x"16d10",-- 5841
x"108c0",-- 4236
x"0ec50",-- 3781
x"16090",-- 5641
x"17c60",-- 6086
x"0f7b0",-- 3963
x"09090",-- 2313
x"088e0",-- 2190
x"070e0",-- 1806
x"04a20",-- 1186
x"04ed0",-- 1261
x"013f0",-- 319
x"f8390",-- -1991
x"f4ed0",-- -2835
x"f8c00",-- -1856
x"f7970",-- -2153
x"f2cd0",-- -3379
x"f35c0",-- -3236
x"f2910",-- -3439
x"ed630",-- -4765
x"edc20",-- -4670
x"f42b0",-- -3029
x"f3e50",-- -3099
x"ef590",-- -4263
x"f06c0",-- -3988
x"f20d0",-- -3571
x"f1040",-- -3836
x"f49b0",-- -2917
x"fa170",-- -1513
x"f7660",-- -2202
x"f3270",-- -3289
x"f7330",-- -2253
x"fc5a0",-- -934
x"fc4b0",-- -949
x"fcf80",-- -776
x"fede0",-- -290
x"fca00",-- -864
x"fb970",-- -1129
x"01cc0",-- 460
x"057b0",-- 1403
x"01db0",-- 475
x"00cb0",-- 203
x"03bd0",-- 957
x"04030",-- 1027
x"03d30",-- 979
x"082f0",-- 2095
x"086e0",-- 2158
x"03bd0",-- 957
x"03260",-- 806
x"080c0",-- 2060
x"06a90",-- 1705
x"04430",-- 1091
x"03e40",-- 996
x"ffc20",-- -62
x"00850",-- 133
x"03a80",-- 936
x"02160",-- 534
x"fb4a0",-- -1206
x"f8d20",-- -1838
x"fa140",-- -1516
x"fb560",-- -1194
x"f92f0",-- -1745
x"f51b0",-- -2789
x"f2370",-- -3529
x"f1de0",-- -3618
x"f31d0",-- -3299
x"f42a0",-- -3030
x"f42b0",-- -3029
x"f1840",-- -3708
x"f1950",-- -3691
x"f5700",-- -2704
x"f7dd0",-- -2083
x"f9d50",-- -1579
x"fcee0",-- -786
x"ff880",-- -120
x"00fc0",-- 252
x"068c0",-- 1676
x"0ab90",-- 2745
x"0d080",-- 3336
x"0f760",-- 3958
x"12c50",-- 4805
x"162c0",-- 5676
x"14ea0",-- 5354
x"17bf0",-- 6079
x"1f1a0",-- 7962
x"21850",-- 8581
x"1be60",-- 7142
x"16fa0",-- 5882
x"1a410",-- 6721
x"1e770",-- 7799
x"1a9a0",-- 6810
x"14b60",-- 5302
x"0ff30",-- 4083
x"0aa90",-- 2729
x"09220",-- 2338
x"0acc0",-- 2764
x"06ea0",-- 1770
x"fcca0",-- -822
x"f7600",-- -2208
x"f8e90",-- -1815
x"f7cb0",-- -2101
x"f4080",-- -3064
x"f2f50",-- -3339
x"f1950",-- -3691
x"ec790",-- -4999
x"eb150",-- -5355
x"ef900",-- -4208
x"f0c30",-- -3901
x"ece80",-- -4888
x"ec350",-- -5067
x"ee050",-- -4603
x"ecfc0",-- -4868
x"edf60",-- -4618
x"f36a0",-- -3222
x"f49e0",-- -2914
x"efca0",-- -4150
x"f0480",-- -4024
x"f5fd0",-- -2563
x"f76a0",-- -2198
x"f76b0",-- -2197
x"fa2a0",-- -1494
x"f9a60",-- -1626
x"f6fc0",-- -2308
x"faeb0",-- -1301
x"016f0",-- 367
x"00410",-- 65
x"fd060",-- -762
x"ff7c0",-- -132
x"01120",-- 274
x"01c90",-- 457
x"02280",-- 552
x"03d30",-- 979
x"05950",-- 1429
x"02f70",-- 759
x"00c50",-- 197
x"01d50",-- 469
x"04230",-- 1059
x"04a40",-- 1188
x"01ea0",-- 490
x"fd4f0",-- -689
x"fc490",-- -951
x"fee80",-- -280
x"00640",-- 100
x"fd200",-- -736
x"f8670",-- -1945
x"f83a0",-- -1990
x"fa480",-- -1464
x"fb620",-- -1182
x"fc460",-- -954
x"fb540",-- -1196
x"fa2a0",-- -1494
x"fca70",-- -857
x"01770",-- 375
x"03900",-- 912
x"04390",-- 1081
x"06c00",-- 1728
x"0af20",-- 2802
x"08a00",-- 2208
x"08a70",-- 2215
x"0cf90",-- 3321
x"14590",-- 5209
x"1afb0",-- 6907
x"17960",-- 6038
x"10cc0",-- 4300
x"10ff0",-- 4351
x"1a0f0",-- 6671
x"20b10",-- 8369
x"1b620",-- 7010
x"0f920",-- 3986
x"0ad90",-- 2777
x"0db00",-- 3504
x"11fb0",-- 4603
x"10000",-- 4096
x"06f90",-- 1785
x"fdda0",-- -550
x"fa1b0",-- -1509
x"fc9e0",-- -866
x"fe370",-- -457
x"fb090",-- -1271
x"f56d0",-- -2707
x"f1650",-- -3739
x"efef0",-- -4113
x"f0f20",-- -3854
x"f4ac0",-- -2900
x"f5220",-- -2782
x"f19d0",-- -3683
x"edd30",-- -4653
x"ee150",-- -4587
x"f14f0",-- -3761
x"f4fd0",-- -2819
x"f6b60",-- -2378
x"f41b0",-- -3045
x"f0b20",-- -3918
x"f10c0",-- -3828
x"f6490",-- -2487
x"fad90",-- -1319
x"fa520",-- -1454
x"f6890",-- -2423
x"f3e70",-- -3097
x"f6700",-- -2448
x"fb9a0",-- -1126
x"ff290",-- -215
x"fccf0",-- -817
x"f8a50",-- -1883
x"f5ae0",-- -2642
x"fc6e0",-- -914
x"ffe90",-- -23
x"fdd60",-- -554
x"fe6b0",-- -405
x"fb950",-- -1131
x"f9920",-- -1646
x"fb2a0",-- -1238
x"fe0a0",-- -502
x"fe9e0",-- -354
x"fea80",-- -344
x"fa660",-- -1434
x"f7400",-- -2240
x"f9110",-- -1775
x"fdfd0",-- -515
x"ffb50",-- -75
x"fbd00",-- -1072
x"f7c40",-- -2108
x"f76b0",-- -2197
x"fd680",-- -664
x"03210",-- 801
x"029b0",-- 667
x"ff110",-- -239
x"ffdb0",-- -37
x"05240",-- 1316
x"0a9d0",-- 2717
x"0eb80",-- 3768
x"0f4f0",-- 3919
x"103c0",-- 4156
x"11f80",-- 4600
x"14110",-- 5137
x"106b0",-- 4203
x"13490",-- 4937
x"22410",-- 8769
x"26e70",-- 9959
x"186d0",-- 6253
x"0d240",-- 3364
x"16fc0",-- 5884
x"26420",-- 9794
x"23fa0",-- 9210
x"14d60",-- 5334
x"0b2b0",-- 2859
x"080c0",-- 2060
x"0bc90",-- 3017
x"11fb0",-- 4603
x"0d9a0",-- 3482
x"fcbb0",-- -837
x"f0820",-- -3966
x"f4de0",-- -2850
x"fb680",-- -1176
x"f7290",-- -2263
x"f0f30",-- -3853
x"ee700",-- -4496
x"e8f30",-- -5901
x"e5d10",-- -6703
x"ed130",-- -4845
x"f3e70",-- -3097
x"eebe0",-- -4418
x"e7060",-- -6394
x"e82d0",-- -6099
x"ec370",-- -5065
x"ee890",-- -4471
x"f3650",-- -3227
x"f5f10",-- -2575
x"efac0",-- -4180
x"e9100",-- -5872
x"ebf90",-- -5127
x"fa210",-- -1503
x"02300",-- 560
x"f9310",-- -1743
x"ec210",-- -5087
x"ebcf0",-- -5169
x"f94a0",-- -1718
x"04870",-- 1159
x"ffe50",-- -27
x"f4f20",-- -2830
x"ef830",-- -4221
x"f5e70",-- -2585
x"01c90",-- 457
x"02b40",-- 692
x"fad20",-- -1326
x"f75b0",-- -2213
x"f6ee0",-- -2322
x"fac60",-- -1338
x"00440",-- 68
x"008f0",-- 143
x"fd240",-- -732
x"fa280",-- -1496
x"fa940",-- -1388
x"fda60",-- -602
x"02f20",-- 754
x"05030",-- 1283
x"014e0",-- 334
x"ff600",-- -160
x"02fc0",-- 764
x"0a820",-- 2690
x"0eb30",-- 3763
x"0f540",-- 3924
x"0e9f0",-- 3743
x"125c0",-- 4700
x"16c70",-- 5831
x"18860",-- 6278
x"17710",-- 6001
x"17270",-- 5927
x"22840",-- 8836
x"28f70",-- 10487
x"21c30",-- 8643
x"18eb0",-- 6379
x"1d370",-- 7479
x"27370",-- 10039
x"28180",-- 10264
x"1c400",-- 7232
x"13620",-- 4962
x"102d0",-- 4141
x"11090",-- 4361
x"12ef0",-- 4847
x"0bea0",-- 3050
x"00410",-- 65
x"f78b0",-- -2165
x"f5ae0",-- -2642
x"f6d00",-- -2352
x"f4260",-- -3034
x"edc90",-- -4663
x"e8b00",-- -5968
x"e6df0",-- -6433
x"e5130",-- -6893
x"e58b0",-- -6773
x"e8730",-- -6029
x"e84c0",-- -6068
x"e3fb0",-- -7173
x"e39a0",-- -7270
x"e6c10",-- -6463
x"e9250",-- -5851
x"ebbf0",-- -5185
x"ee190",-- -4583
x"ecd20",-- -4910
x"e96d0",-- -5779
x"edfe0",-- -4610
x"f5720",-- -2702
x"f5570",-- -2729
x"f1c20",-- -3646
x"f2000",-- -3584
x"f3c50",-- -3131
x"f5840",-- -2684
x"f7680",-- -2200
x"f8930",-- -1901
x"f70e0",-- -2290
x"f5c00",-- -2624
x"f5df0",-- -2593
x"f9040",-- -1788
x"fa200",-- -1504
x"f8a20",-- -1886
x"f9700",-- -1680
x"fa0f0",-- -1521
x"f9ec0",-- -1556
x"fb6f0",-- -1169
x"fcb90",-- -839
x"fe0d0",-- -499
x"fecb0",-- -309
x"ff2e0",-- -210
x"00700",-- 112
x"01e50",-- 485
x"04ae0",-- 1198
x"08c00",-- 2240
x"092c0",-- 2348
x"0a0a0",-- 2570
x"0d4e0",-- 3406
x"12a40",-- 4772
x"15650",-- 5477
x"1af20",-- 6898
x"1ac70",-- 6855
x"15eb0",-- 5611
x"17490",-- 5961
x"1ddf0",-- 7647
x"2baf0",-- 11183
x"2ce70",-- 11495
x"20190",-- 8217
x"19740",-- 6516
x"23030",-- 8963
x"2d3c0",-- 11580
x"2cae0",-- 11438
x"1f240",-- 7972
x"14230",-- 5155
x"11dc0",-- 4572
x"14b40",-- 5300
x"16250",-- 5669
x"0e8c0",-- 3724
x"011f0",-- 287
x"f7060",-- -2298
x"f4930",-- -2925
x"f58e0",-- -2674
x"f3bb0",-- -3141
x"ee780",-- -4488
x"e71b0",-- -6373
x"e1cf0",-- -7729
x"df810",-- -8319
x"e2d80",-- -7464
x"e7db0",-- -6181
x"e5950",-- -6763
x"debf0",-- -8513
x"dca00",-- -9056
x"e0470",-- -8121
x"e6280",-- -6616
x"ea2e0",-- -5586
x"e6c90",-- -6455
x"e4140",-- -7148
x"e4580",-- -7080
x"ead90",-- -5415
x"f1ef0",-- -3601
x"f0b20",-- -3918
x"ed660",-- -4762
x"ed630",-- -4765
x"ef400",-- -4288
x"f50b0",-- -2805
x"f83a0",-- -1990
x"f50e0",-- -2802
x"f2df0",-- -3361
x"f2de0",-- -3362
x"f69b0",-- -2405
x"fba10",-- -1119
x"fb9e0",-- -1122
x"f8e80",-- -1816
x"f7c40",-- -2108
x"fa7a0",-- -1414
x"fefd0",-- -259
x"01b70",-- 439
x"01090",-- 265
x"fef00",-- -272
x"00480",-- 72
x"056f0",-- 1391
x"0a320",-- 2610
x"0c140",-- 3092
x"0a8e0",-- 2702
x"0bb80",-- 3000
x"11210",-- 4385
x"17920",-- 6034
x"1b5f0",-- 7007
x"1e7a0",-- 7802
x"1dba0",-- 7610
x"1a220",-- 6690
x"19f10",-- 6641
x"22b50",-- 8885
x"32830",-- 12931
x"31940",-- 12692
x"21880",-- 8584
x"1ae30",-- 6883
x"25e70",-- 9703
x"32a10",-- 12961
x"2fc10",-- 12225
x"1fc90",-- 8137
x"144b0",-- 5195
x"10f20",-- 4338
x"140c0",-- 5132
x"17e20",-- 6114
x"10570",-- 4183
x"fe8a0",-- -374
x"f1b30",-- -3661
x"f1650",-- -3739
x"f4e90",-- -2839
x"f2e90",-- -3351
x"ec8f0",-- -4977
x"e2e20",-- -7454
x"dbaf0",-- -9297
x"dbf70",-- -9225
x"e2eb0",-- -7445
x"e7e20",-- -6174
x"e2140",-- -7660
x"d9500",-- -9904
x"d9160",-- -9962
x"df4b0",-- -8373
x"e6470",-- -6585
x"e65a0",-- -6566
x"e52a0",-- -6870
x"e18b0",-- -7797
x"df460",-- -8378
x"e9a20",-- -5726
x"f2750",-- -3467
x"efae0",-- -4178
x"e96d0",-- -5779
x"e8da0",-- -5926
x"edd10",-- -4655
x"f5b60",-- -2634
x"f72f0",-- -2257
x"f1e20",-- -3614
x"ee610",-- -4511
x"f2640",-- -3484
x"f8840",-- -1916
x"fc520",-- -942
x"fb420",-- -1214
x"f6d00",-- -2352
x"f82b0",-- -2005
x"fe170",-- -489
x"02ef0",-- 751
x"03e40",-- 996
x"02b20",-- 690
x"02530",-- 595
x"04eb0",-- 1259
x"09ef0",-- 2543
x"0ff30",-- 4083
x"0ffa0",-- 4090
x"0e2c0",-- 3628
x"11450",-- 4421
x"166d0",-- 5741
x"1b880",-- 7048
x"21830",-- 8579
x"22f20",-- 8946
x"1c0f0",-- 7183
x"17c90",-- 6089
x"1f1e0",-- 7966
x"33670",-- 13159
x"38770",-- 14455
x"263b0",-- 9787
x"19760",-- 6518
x"243e0",-- 9278
x"33b10",-- 13233
x"34b50",-- 13493
x"25880",-- 9608
x"17600",-- 5984
x"12140",-- 4628
x"14280",-- 5160
x"18680",-- 6248
x"143e0",-- 5182
x"05180",-- 1304
x"f4940",-- -2924
x"eff10",-- -4111
x"f3d60",-- -3114
x"f3700",-- -3216
x"ee2b0",-- -4565
x"e5d90",-- -6695
x"dbf60",-- -9226
x"d8260",-- -10202
x"de240",-- -8668
x"e6ec0",-- -6420
x"e2e90",-- -7447
x"d8c90",-- -10039
x"d51b0",-- -10981
x"da580",-- -9640
x"e0300",-- -8144
x"e4000",-- -7168
x"e30c0",-- -7412
x"de260",-- -8666
x"dec40",-- -8508
x"e3e80",-- -7192
x"e9200",-- -5856
x"ed150",-- -4843
x"ebdb0",-- -5157
x"e80b0",-- -6133
x"e8c90",-- -5943
x"ed400",-- -4800
x"f1740",-- -3724
x"f4c50",-- -2875
x"f3270",-- -3289
x"ef4a0",-- -4278
x"f14f0",-- -3761
x"f9d80",-- -1576
x"fe0c0",-- -500
x"fcdc0",-- -804
x"fa750",-- -1419
x"fb6d0",-- -1171
x"01680",-- 360
x"06e80",-- 1768
x"09490",-- 2377
x"06ff0",-- 1791
x"06ac0",-- 1708
x"0bc90",-- 3017
x"10e00",-- 4320
x"12f90",-- 4857
x"14ae0",-- 5294
x"15da0",-- 5594
x"18a90",-- 6313
x"1b550",-- 6997
x"22950",-- 8853
x"23d50",-- 9173
x"211a0",-- 8474
x"1d6f0",-- 7535
x"21710",-- 8561
x"313f0",-- 12607
x"36040",-- 13828
x"2a6b0",-- 10859
x"20ed0",-- 8429
x"27580",-- 10072
x"31980",-- 12696
x"32810",-- 12929
x"25060",-- 9478
x"1aa40",-- 6820
x"162f0",-- 5679
x"14c70",-- 5319
x"15880",-- 5512
x"10730",-- 4211
x"03b20",-- 946
x"f6690",-- -2455
x"f1f90",-- -3591
x"f1950",-- -3691
x"eef00",-- -4368
x"eada0",-- -5414
x"e3ac0",-- -7252
x"dc6e0",-- -9106
x"d9040",-- -9980
x"dc100",-- -9200
x"e0bf0",-- -8001
x"df270",-- -8409
x"d83a0",-- -10182
x"d65f0",-- -10657
x"d7d90",-- -10279
x"db640",-- -9372
x"dfde0",-- -8226
x"e21f0",-- -7649
x"e1410",-- -7871
x"ddd90",-- -8743
x"dd520",-- -8878
x"e5750",-- -6795
x"eeed0",-- -4371
x"ec230",-- -5085
x"e5b10",-- -6735
x"e3320",-- -7374
x"e8de0",-- -5922
x"f3a10",-- -3167
x"f6c80",-- -2360
x"efe20",-- -4126
x"ebfe0",-- -5122
x"f0fa0",-- -3846
x"fa7f0",-- -1409
x"00410",-- 65
x"fd970",-- -617
x"f92a0",-- -1750
x"fcd00",-- -816
x"044b0",-- 1099
x"0a110",-- 2577
x"0b2e0",-- 2862
x"09650",-- 2405
x"09450",-- 2373
x"0f100",-- 3856
x"138d0",-- 5005
x"16fe0",-- 5886
x"18250",-- 6181
x"189d0",-- 6301
x"1a890",-- 6793
x"1f7d0",-- 8061
x"26100",-- 9744
x"24750",-- 9333
x"20200",-- 8224
x"1d9b0",-- 7579
x"29a50",-- 10661
x"378a0",-- 14218
x"31d00",-- 12752
x"244f0",-- 9295
x"22ea0",-- 8938
x"2ed80",-- 11992
x"327f0",-- 12927
x"251e0",-- 9502
x"246d0",-- 9325
x"23c80",-- 9160
x"13040",-- 4868
x"0b5d0",-- 2909
x"116f0",-- 4463
x"11c60",-- 4550
x"04710",-- 1137
x"f1510",-- -3759
x"ec1f0",-- -5089
x"eccf0",-- -4913
x"ee210",-- -4575
x"ec8e0",-- -4978
x"e24c0",-- -7604
x"d82b0",-- -10197
x"d4180",-- -11240
x"dd0c0",-- -8948
x"e38b0",-- -7285
x"de8f0",-- -8561
x"d7130",-- -10477
x"d2790",-- -11655
x"d6fb0",-- -10501
x"de7e0",-- -8578
x"e57c0",-- -6788
x"e4880",-- -7032
x"db570",-- -9385
x"d8d70",-- -10025
x"e19d0",-- -7779
x"ee320",-- -4558
x"f11a0",-- -3814
x"e5ab0",-- -6741
x"dd2f0",-- -8913
x"e6dc0",-- -6436
x"f2bb0",-- -3397
x"f5ac0",-- -2644
x"f1f70",-- -3593
x"eca30",-- -4957
x"eaee0",-- -5394
x"f65c0",-- -2468
x"022b0",-- 555
x"ff110",-- -239
x"f9330",-- -1741
x"fa710",-- -1423
x"00d50",-- 213
x"085e0",-- 2142
x"0cf00",-- 3312
x"0bf40",-- 3060
x"072b0",-- 1835
x"0a590",-- 2649
x"13a10",-- 5025
x"17650",-- 5989
x"18340",-- 6196
x"17920",-- 6034
x"19780",-- 6520
x"1c0f0",-- 7183
x"25800",-- 9600
x"27d50",-- 10197
x"21780",-- 8568
x"1e280",-- 7720
x"22110",-- 8721
x"31930",-- 12691
x"37c60",-- 14278
x"2b1a0",-- 11034
x"21ff0",-- 8703
x"27aa0",-- 10154
x"30c50",-- 12485
x"33e90",-- 13289
x"26db0",-- 9947
x"1a7c0",-- 6780
x"15f00",-- 5616
x"16900",-- 5776
x"15fb0",-- 5627
x"0de40",-- 3556
x"03d50",-- 981
x"f7f10",-- -2063
x"f1540",-- -3756
x"f1040",-- -3836
x"ed390",-- -4807
x"e93e0",-- -5826
x"e1d80",-- -7720
x"db900",-- -9328
x"d8800",-- -10112
x"d9d90",-- -9767
x"de440",-- -8636
x"dd040",-- -8956
x"d6080",-- -10744
x"d1630",-- -11933
x"d5110",-- -10991
x"de300",-- -8656
x"e32a0",-- -7382
x"dd700",-- -8848
x"d7e50",-- -10267
x"db4b0",-- -9397
x"e46e0",-- -7058
x"ea870",-- -5497
x"ea760",-- -5514
x"e1d80",-- -7720
x"e0190",-- -8167
x"e9810",-- -5759
x"f1b30",-- -3661
x"f1b60",-- -3658
x"ede20",-- -4638
x"eb180",-- -5352
x"ef540",-- -4268
x"f8e40",-- -1820
x"fe690",-- -407
x"fc050",-- -1019
x"f97a0",-- -1670
x"fc1c0",-- -996
x"036d0",-- 877
x"0a0d0",-- 2573
x"0b920",-- 2962
x"09380",-- 2360
x"09360",-- 2358
x"0e4b0",-- 3659
x"156c0",-- 5484
x"16f40",-- 5876
x"16d10",-- 5841
x"17ce0",-- 6094
x"1b6f0",-- 7023
x"1f870",-- 8071
x"24f60",-- 9462
x"26480",-- 9800
x"226d0",-- 8813
x"1f0b0",-- 7947
x"21df0",-- 8671
x"2fd50",-- 12245
x"37af0",-- 14255
x"2d440",-- 11588
x"21550",-- 8533
x"25d50",-- 9685
x"2fb40",-- 12212
x"357f0",-- 13695
x"29740",-- 10612
x"1af60",-- 6902
x"15530",-- 5459
x"15a50",-- 5541
x"172c0",-- 5932
x"112c0",-- 4396
x"04f50",-- 1269
x"f8760",-- -1930
x"f13d0",-- -3779
x"f1390",-- -3783
x"ef2f0",-- -4305
x"eb450",-- -5307
x"e2fd0",-- -7427
x"d9e10",-- -9759
x"d8010",-- -10239
x"db2a0",-- -9430
x"df200",-- -8416
x"dd640",-- -8860
x"d4c90",-- -11063
x"ce3f0",-- -12737
x"d4220",-- -11230
x"e1830",-- -7805
x"e4a00",-- -7008
x"da1f0",-- -9697
x"d4510",-- -11183
x"da100",-- -9712
x"e7a40",-- -6236
x"ec850",-- -4987
x"e71f0",-- -6369
x"dea80",-- -8536
x"dee20",-- -8478
x"eb590",-- -5287
x"f3a90",-- -3159
x"f1270",-- -3801
x"eb6f0",-- -5265
x"ea440",-- -5564
x"f05c0",-- -4004
x"fa490",-- -1463
x"ff9c0",-- -100
x"fbbd0",-- -1091
x"f87f0",-- -1921
x"fcb40",-- -844
x"049d0",-- 1181
x"0bcc0",-- 3020
x"0ca00",-- 3232
x"08960",-- 2198
x"08b60",-- 2230
x"0f4a0",-- 3914
x"163e0",-- 5694
x"18720",-- 6258
x"16e60",-- 5862
x"173c0",-- 5948
x"1c9a0",-- 7322
x"201d0",-- 8221
x"24f20",-- 9458
x"25c10",-- 9665
x"22790",-- 8825
x"1ec90",-- 7881
x"23210",-- 8993
x"2f690",-- 12137
x"36920",-- 13970
x"2cc20",-- 11458
x"21e10",-- 8673
x"26400",-- 9792
x"2f7a0",-- 12154
x"33f30",-- 13299
x"28520",-- 10322
x"1acf0",-- 6863
x"151f0",-- 5407
x"158d0",-- 5517
x"16950",-- 5781
x"10020",-- 4098
x"03a80",-- 936
x"f80c0",-- -2036
x"f19f0",-- -3681
x"f1240",-- -3804
x"eea70",-- -4441
x"e9ef0",-- -5649
x"e2a30",-- -7517
x"d9f70",-- -9737
x"d7ca0",-- -10294
x"db2f0",-- -9425
x"de530",-- -8621
x"dbc70",-- -9273
x"cf230",-- -12509
x"cf9a0",-- -12390
x"de410",-- -8639
x"e0600",-- -8096
x"d9e80",-- -9752
x"d7430",-- -10429
x"d7390",-- -10439
x"e00b0",-- -8181
x"eaa50",-- -5467
x"e5090",-- -6903
x"dd770",-- -8841
x"e0ad0",-- -8019
x"e85a0",-- -6054
x"ee580",-- -4520
x"efe70",-- -4121
x"ec7d0",-- -4995
x"e9ca0",-- -5686
x"efab0",-- -4181
x"f87a0",-- -1926
x"fb9c0",-- -1124
x"fad70",-- -1321
x"fa7d0",-- -1411
x"fd4e0",-- -690
x"014c0",-- 332
x"07b70",-- 1975
x"0c730",-- 3187
x"08930",-- 2195
x"073f0",-- 1855
x"0e1b0",-- 3611
x"14090",-- 5129
x"14ac0",-- 5292
x"15dd0",-- 5597
x"160a0",-- 5642
x"19300",-- 6448
x"1faa0",-- 8106
x"22650",-- 8805
x"237e0",-- 9086
x"1fa00",-- 8096
x"203b0",-- 8251
x"23010",-- 8961
x"27800",-- 10112
x"2e6b0",-- 11883
x"30840",-- 12420
x"27150",-- 10005
x"22d90",-- 8921
x"2a720",-- 10866
x"318c0",-- 12684
x"2db40",-- 11700
x"21620",-- 8546
x"18e30",-- 6371
x"15440",-- 5444
x"16f40",-- 5876
x"16090",-- 5641
x"0ab60",-- 2742
x"fd880",-- -632
x"f6190",-- -2535
x"f32c0",-- -3284
x"f1f40",-- -3596
x"ee2b0",-- -4565
x"e6b90",-- -6471
x"de0f0",-- -8689
x"da580",-- -9640
x"db4b0",-- -9397
x"de3f0",-- -8641
x"dc4c0",-- -9140
x"d38b0",-- -11381
x"d1000",-- -12032
x"dae70",-- -9497
x"def80",-- -8456
x"da920",-- -9582
x"d79f0",-- -10337
x"d8a30",-- -10077
x"df160",-- -8426
x"e5f40",-- -6668
x"e4330",-- -7117
x"deee0",-- -8466
x"e26f0",-- -7569
x"e8990",-- -5991
x"e97f0",-- -5761
x"ecd50",-- -4907
x"ee980",-- -4456
x"ec8e0",-- -4978
x"ef250",-- -4315
x"f4bc0",-- -2884
x"f8050",-- -2043
x"fac30",-- -1341
x"fd060",-- -762
x"fd630",-- -669
x"fed20",-- -302
x"041c0",-- 1052
x"09e50",-- 2533
x"09d10",-- 2513
x"08f90",-- 2297
x"0b3b0",-- 2875
x"10400",-- 4160
x"13a30",-- 5027
x"142c0",-- 5164
x"16950",-- 5781
x"182c0",-- 6188
x"1bc90",-- 7113
x"1f010",-- 7937
x"22ca0",-- 8906
x"22110",-- 8721
x"1e980",-- 7832
x"21830",-- 8579
x"24930",-- 9363
x"29880",-- 10632
x"2f0f0",-- 12047
x"2ab60",-- 10934
x"24810",-- 9345
x"26e70",-- 9959
x"2cbb0",-- 11451
x"2ef40",-- 12020
x"27290",-- 10025
x"1e110",-- 7697
x"176a0",-- 5994
x"162d0",-- 5677
x"17aa0",-- 6058
x"10ed0",-- 4333
x"04940",-- 1172
x"faf30",-- -1293
x"f5ec0",-- -2580
x"f41b0",-- -3045
x"f0d70",-- -3881
x"ebdd0",-- -5155
x"e2af0",-- -7505
x"dd550",-- -8875
x"dca00",-- -9056
x"de210",-- -8671
x"ddb30",-- -8781
x"d65f0",-- -10657
x"d4f10",-- -11023
x"da6e0",-- -9618
x"dc2d0",-- -9171
x"d9f90",-- -9735
x"d9ca0",-- -9782
x"da920",-- -9582
x"de100",-- -8688
x"e2530",-- -7597
x"e23f0",-- -7617
x"dfcc0",-- -8244
x"e2e60",-- -7450
x"e73b0",-- -6341
x"e8640",-- -6044
x"ea4c0",-- -5556
x"ec600",-- -5024
x"ec740",-- -5004
x"eeb20",-- -4430
x"f2bc0",-- -3396
x"f60c0",-- -2548
x"f8210",-- -2015
x"faca0",-- -1334
x"fcc00",-- -832
x"febb0",-- -325
x"02b10",-- 689
x"06d20",-- 1746
x"07da0",-- 2010
x"08b60",-- 2230
x"0c1e0",-- 3102
x"0ecf0",-- 3791
x"11df0",-- 4575
x"13150",-- 4885
x"14f90",-- 5369
x"18280",-- 6184
x"1c090",-- 7177
x"1de70",-- 7655
x"1eba0",-- 7866
x"21560",-- 8534
x"21b90",-- 8633
x"21ba0",-- 8634
x"22cc0",-- 8908
x"25dc0",-- 9692
x"2bf80",-- 11256
x"2da30",-- 11683
x"27370",-- 10039
x"24ed0",-- 9453
x"29410",-- 10561
x"2d9d0",-- 11677
x"2a770",-- 10871
x"204b0",-- 8267
x"19670",-- 6503
x"172b0",-- 5931
x"16c00",-- 5824
x"13080",-- 4872
x"08a40",-- 2212
x"fdd50",-- -555
x"f7560",-- -2218
x"f5b60",-- -2634
x"f2e30",-- -3357
x"ebe80",-- -5144
x"e5160",-- -6890
x"e0080",-- -8184
x"de5d0",-- -8611
x"ddd10",-- -8751
x"dcb20",-- -9038
x"d8ab0",-- -10069
x"d6da0",-- -10534
x"d8ad0",-- -10067
x"db0c0",-- -9460
x"db900",-- -9328
x"d9750",-- -9867
x"da2e0",-- -9682
x"dd6d0",-- -8851
x"df7c0",-- -8324
x"e26e0",-- -7570
x"e2550",-- -7595
x"e0790",-- -8071
x"e5190",-- -6887
x"e8e80",-- -5912
x"e8e80",-- -5912
x"ebac0",-- -5204
x"ed4d0",-- -4787
x"ecc50",-- -4923
x"f0940",-- -3948
x"f5f60",-- -2570
x"f7660",-- -2202
x"f9810",-- -1663
x"fc800",-- -896
x"fe0c0",-- -500
x"01a30",-- 419
x"053f0",-- 1343
x"077b0",-- 1915
x"095e0",-- 2398
x"0ad70",-- 2775
x"0d2c0",-- 3372
x"10de0",-- 4318
x"13120",-- 4882
x"137b0",-- 4987
x"162c0",-- 5676
x"19ab0",-- 6571
x"1c910",-- 7313
x"1e700",-- 7792
x"218a0",-- 8586
x"20520",-- 8274
x"1ea20",-- 7842
x"20fe0",-- 8446
x"24db0",-- 9435
x"2a9f0",-- 10911
x"2c9f0",-- 11423
x"25f30",-- 9715
x"21e40",-- 8676
x"27c90",-- 10185
x"2e450",-- 11845
x"2ba20",-- 11170
x"21100",-- 8464
x"19600",-- 6496
x"17320",-- 5938
x"18320",-- 6194
x"15640",-- 5476
x"0c0f0",-- 3087
x"ffa30",-- -93
x"f8c30",-- -1853
x"f7510",-- -2223
x"f4e90",-- -2839
x"ee760",-- -4490
x"e7e20",-- -6174
x"e19d0",-- -7779
x"de6a0",-- -8598
x"dec10",-- -8511
x"de5b0",-- -8613
x"dc060",-- -9210
x"d8b40",-- -10060
x"d8260",-- -10202
x"d8820",-- -10110
x"dc1f0",-- -9185
x"ddd30",-- -8749
x"dbc00",-- -9280
x"db140",-- -9452
x"de670",-- -8601
x"e1050",-- -7931
x"e44e0",-- -7090
x"e5630",-- -6813
x"e35e0",-- -7330
x"e4fa0",-- -6918
x"e8f30",-- -5901
x"ec6e0",-- -5010
x"ee440",-- -4540
x"ee2d0",-- -4563
x"eeb20",-- -4430
x"f20b0",-- -3573
x"f6d40",-- -2348
x"fa910",-- -1391
x"fc520",-- -942
x"fca30",-- -861
x"fe9b0",-- -357
x"03620",-- 866
x"077b0",-- 1915
x"09150",-- 2325
x"0a070",-- 2567
x"0aed0",-- 2797
x"0dc60",-- 3526
x"122a0",-- 4650
x"14860",-- 5254
x"15880",-- 5512
x"16130",-- 5651
x"1acd0",-- 6861
x"1d240",-- 7460
x"207e0",-- 8318
x"21620",-- 8546
x"1d330",-- 7475
x"1f490",-- 8009
x"255f0",-- 9567
x"270d0",-- 9997
x"2a200",-- 10784
x"289a0",-- 10394
x"24a90",-- 9385
x"26520",-- 9810
x"29c30",-- 10691
x"2b7d0",-- 11133
x"25330",-- 9523
x"1d4e0",-- 7502
x"17ff0",-- 6143
x"16a50",-- 5797
x"16220",-- 5666
x"0f1c0",-- 3868
x"04bb0",-- 1211
x"fc020",-- -1022
x"f6fc0",-- -2308
x"f67b0",-- -2437
x"f1470",-- -3769
x"ea490",-- -5559
x"e4c60",-- -6970
x"e0370",-- -8137
x"df630",-- -8349
x"dfbb0",-- -8261
x"dd180",-- -8936
x"da240",-- -9692
x"da2d0",-- -9683
x"d9900",-- -9840
x"d8fd0",-- -9987
x"dd780",-- -8840
x"df9c0",-- -8292
x"dbfb0",-- -9221
x"db840",-- -9340
x"e0780",-- -8072
x"e3a70",-- -7257
x"e4240",-- -7132
x"e5e80",-- -6680
x"e4260",-- -7130
x"e5810",-- -6783
x"ec440",-- -5052
x"ee640",-- -4508
x"eca50",-- -4955
x"edce0",-- -4658
x"f1f20",-- -3598
x"f4c80",-- -2872
x"f8530",-- -1965
x"fb450",-- -1211
x"fbfd0",-- -1027
x"fe2b0",-- -469
x"01d00",-- 464
x"05c70",-- 1479
x"08bb0",-- 2235
x"09ad0",-- 2477
x"0a210",-- 2593
x"0c7f0",-- 3199
x"11290",-- 4393
x"157e0",-- 5502
x"15470",-- 5447
x"14c30",-- 5315
x"19560",-- 6486
x"1db40",-- 7604
x"20790",-- 8313
x"1f3f0",-- 7999
x"1c810",-- 7297
x"20520",-- 8274
x"25210",-- 9505
x"25f60",-- 9718
x"28790",-- 10361
x"27510",-- 10065
x"252e0",-- 9518
x"27b20",-- 10162
x"28fc0",-- 10492
x"28fe0",-- 10494
x"251c0",-- 9500
x"1fbc0",-- 8124
x"1a1d0",-- 6685
x"16ca0",-- 5834
x"15a10",-- 5537
x"102f0",-- 4143
x"07120",-- 1810
x"fe4e0",-- -434
x"f8110",-- -2031
x"f66e0",-- -2450
x"f37e0",-- -3202
x"ec300",-- -5072
x"e5ae0",-- -6738
x"e1880",-- -7800
x"e0730",-- -8077
x"e0e10",-- -7967
x"de6f0",-- -8593
x"dac30",-- -9533
x"d9700",-- -9872
x"dab20",-- -9550
x"db250",-- -9435
x"dcad0",-- -9043
x"de290",-- -8663
x"dcff0",-- -8961
x"dbaa0",-- -9302
x"df1b0",-- -8421
x"e4880",-- -7032
x"e4a50",-- -7003
x"e4a50",-- -7003
x"e4d00",-- -6960
x"e54a0",-- -6838
x"eb390",-- -5319
x"ef290",-- -4311
x"ed700",-- -4752
x"ed2f0",-- -4817
x"f0480",-- -4024
x"f5160",-- -2794
x"f9070",-- -1785
x"fb3e0",-- -1218
x"fbb30",-- -1101
x"fd060",-- -762
x"01f60",-- 502
x"06580",-- 1624
x"07da0",-- 2010
x"08e60",-- 2278
x"0aef0",-- 2799
x"0dc60",-- 3526
x"10040",-- 4100
x"138a0",-- 5002
x"15a50",-- 5541
x"16af0",-- 5807
x"18a00",-- 6304
x"1b560",-- 6998
x"208e0",-- 8334
x"20720",-- 8306
x"1b910",-- 7057
x"1ec40",-- 7876
x"25500",-- 9552
x"25f30",-- 9715
x"273f0",-- 10047
x"26b80",-- 9912
x"23ff0",-- 9215
x"26f90",-- 9977
x"29c50",-- 10693
x"28f60",-- 10486
x"24070",-- 9223
x"1dbf0",-- 7615
x"19aa0",-- 6570
x"18a90",-- 6313
x"16140",-- 5652
x"0eb60",-- 3766
x"06480",-- 1608
x"ff6f0",-- -145
x"f9900",-- -1648
x"f6f30",-- -2317
x"f3900",-- -3184
x"ed2c0",-- -4820
x"e7150",-- -6379
x"e21a0",-- -7654
x"e1e70",-- -7705
x"e2190",-- -7655
x"dec80",-- -8504
x"dbcf0",-- -9265
x"dc970",-- -9065
x"d93e0",-- -9922
x"d9160",-- -9962
x"e0e90",-- -7959
x"e0150",-- -8171
x"dbe50",-- -9243
x"de1e0",-- -8674
x"dc910",-- -9071
x"e1f20",-- -7694
x"eb630",-- -5277
x"e71f0",-- -6369
x"e05a0",-- -8102
x"e49c0",-- -7012
x"ebce0",-- -5170
x"ef830",-- -4221
x"f1540",-- -3756
x"ed590",-- -4775
x"ec140",-- -5100
x"f44d0",-- -2995
x"fb240",-- -1244
x"fcfc0",-- -772
x"fc4e0",-- -946
x"fabc0",-- -1348
x"ff540",-- -172
x"06f50",-- 1781
x"09a10",-- 2465
x"093f0",-- 2367
x"09220",-- 2338
x"0a210",-- 2593
x"0ee30",-- 3811
x"15620",-- 5474
x"16690",-- 5737
x"149f0",-- 5279
x"16d90",-- 5849
x"19240",-- 6436
x"20a20",-- 8354
x"21c40",-- 8644
x"1a630",-- 6755
x"1c980",-- 7320
x"23bf0",-- 9151
x"265b0",-- 9819
x"28c00",-- 10432
x"25670",-- 9575
x"22460",-- 8774
x"276f0",-- 10095
x"296e0",-- 10606
x"28860",-- 10374
x"22d90",-- 8921
x"1d2b0",-- 7467
x"1a690",-- 6761
x"18cc0",-- 6348
x"148e0",-- 5262
x"0d710",-- 3441
x"07bf0",-- 1983
x"ffdf0",-- -33
x"f8a30",-- -1885
x"f79c0",-- -2148
x"f3390",-- -3271
x"ec4c0",-- -5044
x"e9220",-- -5854
x"e43f0",-- -7105
x"e0d80",-- -7976
x"e1dd0",-- -7715
x"e2490",-- -7607
x"dcc10",-- -9023
x"d8240",-- -10204
x"dc730",-- -9101
x"dfe30",-- -8221
x"df000",-- -8448
x"ddaa0",-- -8790
x"dc260",-- -9178
x"de170",-- -8681
x"e3b30",-- -7245
x"e5d60",-- -6698
x"e26e0",-- -7570
x"e2c90",-- -7479
x"e6ff0",-- -6401
x"e93d0",-- -5827
x"ec580",-- -5032
x"ed630",-- -4765
x"eb4a0",-- -5302
x"ef8b0",-- -4213
x"f3360",-- -3274
x"f5020",-- -2814
x"f8070",-- -2041
x"f9db0",-- -1573
x"fb650",-- -1179
x"fe3c0",-- -452
x"02b10",-- 689
x"04430",-- 1091
x"06870",-- 1671
x"09560",-- 2390
x"091f0",-- 2335
x"0ca70",-- 3239
x"10750",-- 4213
x"12460",-- 4678
x"14180",-- 5144
x"14e30",-- 5347
x"17f50",-- 6133
x"1bc30",-- 7107
x"21820",-- 8578
x"1d000",-- 7424
x"173c0",-- 5948
x"20bd0",-- 8381
x"278d0",-- 10125
x"25830",-- 9603
x"25510",-- 9553
x"22600",-- 8800
x"237e0",-- 9086
x"29960",-- 10646
x"29ca0",-- 10698
x"25ec0",-- 9708
x"1f670",-- 8039
x"1d2e0",-- 7470
x"1a950",-- 6805
x"178c0",-- 6028
x"14e00",-- 5344
x"0d270",-- 3367
x"039e0",-- 926
x"fdc40",-- -572
x"fb3e0",-- -1218
x"f8120",-- -2030
x"f1e70",-- -3609
x"ec8c0",-- -4980
x"e6e90",-- -6423
x"e3540",-- -7340
x"e43c0",-- -7108
x"e3e20",-- -7198
x"e0ab0",-- -8021
x"dcaa0",-- -9046
x"dac30",-- -9533
x"d9140",-- -9964
x"de370",-- -8649
x"e61a0",-- -6630
x"df2d0",-- -8403
x"d9640",-- -9884
x"ddc70",-- -8761
x"e1020",-- -7934
x"e88d0",-- -6003
x"eb310",-- -5327
x"e2470",-- -7609
x"de5f0",-- -8609
x"e8530",-- -6061
x"f1950",-- -3691
x"efcf0",-- -4145
x"ed6d0",-- -4755
x"ec890",-- -4983
x"ee420",-- -4542
x"f7c70",-- -2105
x"fcb10",-- -847
x"fb600",-- -1184
x"f98d0",-- -1651
x"faf20",-- -1294
x"02930",-- 659
x"08870",-- 2183
x"09300",-- 2352
x"071c0",-- 1820
x"078d0",-- 1933
x"0b6c0",-- 2924
x"10860",-- 4230
x"16730",-- 5747
x"13cd0",-- 5069
x"125f0",-- 4703
x"169d0",-- 5789
x"1d580",-- 7512
x"22520",-- 8786
x"1b210",-- 6945
x"18d40",-- 6356
x"21870",-- 8583
x"24810",-- 9345
x"25b20",-- 9650
x"262f0",-- 9775
x"21f80",-- 8696
x"24890",-- 9353
x"28100",-- 10256
x"27eb0",-- 10219
x"23d50",-- 9173
x"1fdd0",-- 8157
x"1bcd0",-- 7117
x"173c0",-- 5948
x"16ea0",-- 5866
x"117e0",-- 4478
x"098a0",-- 2442
x"03fb0",-- 1019
x"fbe00",-- -1056
x"f8760",-- -1930
x"f6b40",-- -2380
x"f0370",-- -4041
x"eaa60",-- -5466
x"e78e0",-- -6258
x"e4e40",-- -6940
x"e23d0",-- -7619
x"e32c0",-- -7380
x"e2000",-- -7680
x"dd040",-- -8956
x"da5a0",-- -9638
x"db870",-- -9337
x"e2670",-- -7577
x"e4460",-- -7098
x"dd070",-- -8953
x"dc0b0",-- -9205
x"dfb10",-- -8271
x"e3ce0",-- -7218
x"ead40",-- -5420
x"e7f40",-- -6156
x"df1e0",-- -8418
x"e39f0",-- -7265
x"eeb70",-- -4425
x"f0550",-- -4011
x"ee240",-- -4572
x"edf20",-- -4622
x"ed840",-- -4732
x"f32c0",-- -3284
x"fb570",-- -1193
x"fb9e0",-- -1122
x"f9340",-- -1740
x"faa70",-- -1369
x"ff7c0",-- -132
x"05f60",-- 1526
x"07fd0",-- 2045
x"06730",-- 1651
x"06f20",-- 1778
x"0aaf0",-- 2735
x"0de70",-- 3559
x"11f80",-- 4600
x"14d70",-- 5335
x"12c50",-- 4805
x"139e0",-- 5022
x"19f10",-- 6641
x"213c0",-- 8508
x"1b060",-- 6918
x"16b90",-- 5817
x"20d30",-- 8403
x"24ac0",-- 9388
x"21ad0",-- 8621
x"24a10",-- 9377
x"23620",-- 9058
x"23ce0",-- 9166
x"28100",-- 10256
x"269f0",-- 9887
x"23d30",-- 9171
x"207c0",-- 8316
x"1f100",-- 7952
x"1a720",-- 6770
x"16980",-- 5784
x"12b30",-- 4787
x"0c700",-- 3184
x"07c70",-- 1991
x"00410",-- 65
x"f90e0",-- -1778
x"f77f0",-- -2177
x"f3f60",-- -3082
x"ee190",-- -4583
x"e8ad0",-- -5971
x"e6000",-- -6656
x"e47b0",-- -7045
x"e3c00",-- -7232
x"e3160",-- -7402
x"de500",-- -8624
x"db410",-- -9407
x"de710",-- -8591
x"e1bb0",-- -7749
x"e0790",-- -8071
x"de460",-- -8634
x"de7b0",-- -8581
x"e1860",-- -7802
x"e3e70",-- -7193
x"e5c40",-- -6716
x"e5fb0",-- -6661
x"e53d0",-- -6851
x"e6050",-- -6651
x"ea620",-- -5534
x"eddd0",-- -4643
x"edc70",-- -4665
x"ee260",-- -4570
x"ef9a0",-- -4198
x"f3130",-- -3309
x"f7720",-- -2190
x"f91d0",-- -1763
x"f98d0",-- -1651
x"fbb30",-- -1101
x"ff710",-- -143
x"022b0",-- 555
x"04170",-- 1047
x"05950",-- 1429
x"07210",-- 1825
x"09c90",-- 2505
x"0c9b0",-- 3227
x"0d030",-- 3331
x"0f770",-- 3959
x"12690",-- 4713
x"15bc0",-- 5564
x"17290",-- 5929
x"1a250",-- 6693
x"1ca20",-- 7330
x"17d70",-- 6103
x"1aec0",-- 6892
x"23300",-- 9008
x"24020",-- 9218
x"21f50",-- 8693
x"22000",-- 8704
x"22520",-- 8786
x"263b0",-- 9787
x"27260",-- 10022
x"26830",-- 9859
x"22790",-- 8825
x"1c840",-- 7300
x"1a520",-- 6738
x"19d80",-- 6616
x"17d00",-- 6096
x"0f060",-- 3846
x"08020",-- 2050
x"02dc0",-- 732
x"fc460",-- -954
x"fa960",-- -1386
x"f8480",-- -1976
x"f0490",-- -4023
x"e8f00",-- -5904
x"e7a20",-- -6238
x"e7bf0",-- -6209
x"e5f60",-- -6666
x"e3ed0",-- -7187
x"e0080",-- -8184
x"dd480",-- -8888
x"de000",-- -8704
x"e11e0",-- -7906
x"e2eb0",-- -7445
x"dfac0",-- -8276
x"ddbb0",-- -8773
x"e1480",-- -7864
x"e3270",-- -7385
x"e5520",-- -6830
x"e79d0",-- -6243
x"e6740",-- -6540
x"e5160",-- -6890
x"e7ac0",-- -6228
x"ed090",-- -4855
x"eedf0",-- -4385
x"ef570",-- -4265
x"efb80",-- -4168
x"efab0",-- -4181
x"f4260",-- -3034
x"f9db0",-- -1573
x"fc350",-- -971
x"fb3b0",-- -1221
x"fad20",-- -1326
x"ff270",-- -217
x"04710",-- 1137
x"076c0",-- 1900
x"07a30",-- 1955
x"065a0",-- 1626
x"08370",-- 2103
x"0ca50",-- 3237
x"126d0",-- 4717
x"138c0",-- 5004
x"11e70",-- 4583
x"135d0",-- 4957
x"190b0",-- 6411
x"1e4f0",-- 7759
x"195f0",-- 6495
x"187f0",-- 6271
x"1fd00",-- 8144
x"22f20",-- 8946
x"23140",-- 8980
x"22630",-- 8803
x"21080",-- 8456
x"251a0",-- 9498
x"27f50",-- 10229
x"26090",-- 9737
x"21010",-- 8449
x"1de40",-- 7652
x"1cd40",-- 7380
x"19f80",-- 6648
x"17af0",-- 6063
x"0fd70",-- 4055
x"08d10",-- 2257
x"05fe0",-- 1534
x"ffea0",-- -22
x"fb250",-- -1243
x"f72c0",-- -2260
x"f1a60",-- -3674
x"ec710",-- -5007
x"e9450",-- -5819
x"e9090",-- -5879
x"e6300",-- -6608
x"e2e90",-- -7447
x"e0870",-- -8057
x"dfb10",-- -8271
x"dfe80",-- -8216
x"e0410",-- -8127
x"e1ba0",-- -7750
x"e0080",-- -8184
x"ddd60",-- -8746
x"e1410",-- -7871
x"e42d0",-- -7123
x"e4880",-- -7032
x"e4940",-- -7020
x"e4ec0",-- -6932
x"e7700",-- -6288
x"e8de0",-- -5922
x"eb040",-- -5372
x"ee210",-- -4575
x"edd60",-- -4650
x"ee8e0",-- -4466
x"f2800",-- -3456
x"f5c40",-- -2620
x"f72a0",-- -2262
x"f9940",-- -1644
x"fb520",-- -1198
x"fc700",-- -912
x"00da0",-- 218
x"04b80",-- 1208
x"04980",-- 1176
x"05bd0",-- 1469
x"084e0",-- 2126
x"0a590",-- 2649
x"0ca50",-- 3237
x"0f9a0",-- 3994
x"11df0",-- 4575
x"13cb0",-- 5067
x"14950",-- 5269
x"16b60",-- 5814
x"1bfd0",-- 7165
x"19550",-- 6485
x"17530",-- 5971
x"1f730",-- 8051
x"24270",-- 9255
x"1fc60",-- 8134
x"1e860",-- 7814
x"22560",-- 8790
x"26450",-- 9797
x"24f60",-- 9462
x"235d0",-- 9053
x"21510",-- 8529
x"1dc10",-- 7617
x"1b910",-- 7057
x"19e20",-- 6626
x"183e0",-- 6206
x"10520",-- 4178
x"07c60",-- 1990
x"06110",-- 1553
x"014f0",-- 335
x"fb310",-- -1231
x"f7f80",-- -2056
x"f2c30",-- -3389
x"ec6a0",-- -5014
x"e9e70",-- -5657
x"ea440",-- -5564
x"e6420",-- -6590
x"e36f0",-- -7313
x"e38d0",-- -7283
x"e07e0",-- -8066
x"df250",-- -8411
x"e0da0",-- -7974
x"e12a0",-- -7894
x"e1880",-- -7800
x"e1220",-- -7902
x"e0290",-- -8151
x"e1e70",-- -7705
x"e4790",-- -7047
x"e67d0",-- -6531
x"e80b0",-- -6133
x"e7510",-- -6319
x"e5c40",-- -6716
x"ea490",-- -5559
x"f0430",-- -4029
x"efed0",-- -4115
x"efdb0",-- -4133
x"f13b0",-- -3781
x"f2ee0",-- -3346
x"f87a0",-- -1926
x"fd950",-- -619
x"fb830",-- -1149
x"fa8c0",-- -1396
x"ff650",-- -155
x"03d10",-- 977
x"06050",-- 1541
x"07360",-- 1846
x"069a0",-- 1690
x"08cc0",-- 2252
x"0c700",-- 3184
x"0ee00",-- 3808
x"120e0",-- 4622
x"13540",-- 4948
x"12840",-- 4740
x"15940",-- 5524
x"1c160",-- 7190
x"18f50",-- 6389
x"16de0",-- 5854
x"1e700",-- 7792
x"221d0",-- 8733
x"21100",-- 8464
x"20040",-- 8196
x"1fc30",-- 8131
x"244c0",-- 9292
x"26ce0",-- 9934
x"24830",-- 9347
x"20520",-- 8274
x"1c8c0",-- 7308
x"1c900",-- 7312
x"1b470",-- 6983
x"178a0",-- 6026
x"106e0",-- 4206
x"09560",-- 2390
x"07210",-- 1825
x"01d80",-- 472
x"fb810",-- -1151
x"f8be0",-- -1858
x"f4710",-- -2959
x"edfe0",-- -4610
x"e9a70",-- -5721
x"e8eb0",-- -5909
x"e76a0",-- -6294
x"e6280",-- -6616
x"e3860",-- -7290
x"deaa0",-- -8534
x"df6b0",-- -8341
x"e1700",-- -7824
x"e1fc0",-- -7684
x"e2b40",-- -7500
x"df610",-- -8351
x"ddd90",-- -8743
x"e3650",-- -7323
x"e7240",-- -6364
x"e6000",-- -6656
x"e3e00",-- -7200
x"e6420",-- -6590
x"e9660",-- -5786
x"ec210",-- -5087
x"efa10",-- -4191
x"eef20",-- -4366
x"ee4e0",-- -4530
x"f32a0",-- -3286
x"f7a40",-- -2140
x"f8f00",-- -1808
x"fa6c0",-- -1428
x"fb480",-- -1208
x"fc530",-- -941
x"00570",-- 87
x"05800",-- 1408
x"06020",-- 1538
x"05e20",-- 1506
x"065d0",-- 1629
x"081c0",-- 2076
x"0cd90",-- 3289
x"11080",-- 4360
x"103c0",-- 4156
x"10900",-- 4240
x"13ba0",-- 5050
x"16eb0",-- 5867
x"1b030",-- 6915
x"184d0",-- 6221
x"16910",-- 5777
x"1ce00",-- 7392
x"22f70",-- 8951
x"21d20",-- 8658
x"1d730",-- 7539
x"1dc40",-- 7620
x"267e0",-- 9854
x"27560",-- 10070
x"222d0",-- 8749
x"1f0a0",-- 7946
x"1cb40",-- 7348
x"1cf40",-- 7412
x"1b5f0",-- 7007
x"16750",-- 5749
x"0e570",-- 3671
x"09f10",-- 2545
x"07180",-- 1816
x"01c90",-- 457
x"fc0c0",-- -1012
x"f73d0",-- -2243
x"f3750",-- -3211
x"ef570",-- -4265
x"ea420",-- -5566
x"e8600",-- -6048
x"e8510",-- -6063
x"e5920",-- -6766
x"e21c0",-- -7652
x"e06a0",-- -8086
x"e0710",-- -8079
x"e1790",-- -7815
x"e3400",-- -7360
x"e1610",-- -7839
x"de1e0",-- -8674
x"e0820",-- -8062
x"e4c90",-- -6967
x"e54c0",-- -6836
x"e4940",-- -7020
x"e5c50",-- -6715
x"e7270",-- -6361
x"e9d90",-- -5671
x"ede80",-- -4632
x"ef130",-- -4333
x"eeed0",-- -4371
x"f0ac0",-- -3924
x"f4910",-- -2927
x"f7f80",-- -2056
x"fa840",-- -1404
x"fabb0",-- -1349
x"fb010",-- -1279
x"ff3a0",-- -198
x"035e0",-- 862
x"03c90",-- 969
x"03f80",-- 1016
x"069f0",-- 1695
x"08fa0",-- 2298
x"0a190",-- 2585
x"0ce60",-- 3302
x"0f620",-- 3938
x"0fc90",-- 4041
x"137e0",-- 4990
x"15350",-- 5429
x"16720",-- 5746
x"18b30",-- 6323
x"171c0",-- 5916
x"18bb0",-- 6331
x"1e040",-- 7684
x"20770",-- 8311
x"220c0",-- 8716
x"1efb0",-- 7931
x"1beb0",-- 7147
x"22f60",-- 8950
x"28570",-- 10327
x"25010",-- 9473
x"1aef0",-- 6895
x"18450",-- 6213
x"1a2a0",-- 6698
x"1a9d0",-- 6813
x"1a230",-- 6691
x"0f950",-- 3989
x"028f0",-- 655
x"ffe90",-- -23
x"01300",-- 304
x"fffe0",-- -2
x"f8e30",-- -1821
x"ef020",-- -4350
x"e91b0",-- -5861
x"e7ef0",-- -6161
x"ec0d0",-- -5107
x"eb150",-- -5355
x"e42b0",-- -7125
x"dded0",-- -8723
x"ddc00",-- -8768
x"e2060",-- -7674
x"e5330",-- -6861
x"e4850",-- -7035
x"df660",-- -8346
x"dd570",-- -8873
x"e1e70",-- -7705
x"e6df0",-- -6433
x"e8050",-- -6139
x"e5890",-- -6775
x"e5400",-- -6848
x"e8080",-- -6136
x"ebec0",-- -5140
x"f1770",-- -3721
x"f2640",-- -3484
x"eff90",-- -4103
x"f0c10",-- -3903
x"f58b0",-- -2677
x"fbdd0",-- -1059
x"fc8a0",-- -886
x"fb650",-- -1179
x"fc260",-- -986
x"fe7d0",-- -387
x"032c0",-- 812
x"06bb0",-- 1723
x"07530",-- 1875
x"05c20",-- 1474
x"06890",-- 1673
x"0b010",-- 2817
x"0e5e0",-- 3678
x"0f650",-- 3941
x"11490",-- 4425
x"12d90",-- 4825
x"12d90",-- 4825
x"16890",-- 5769
x"18700",-- 6256
x"173c0",-- 5948
x"1bfd0",-- 7165
x"1e820",-- 7810
x"1b6c0",-- 7020
x"1ce20",-- 7394
x"20cc0",-- 8396
x"23670",-- 9063
x"23ab0",-- 9131
x"20c40",-- 8388
x"20660",-- 8294
x"1d1f0",-- 7455
x"1bdd0",-- 7133
x"1af10",-- 6897
x"16910",-- 5777
x"11830",-- 4483
x"0b950",-- 2965
x"069b0",-- 1691
x"04890",-- 1161
x"00ca0",-- 202
x"f9a90",-- -1623
x"f34f0",-- -3249
x"f17f0",-- -3713
x"ed8e0",-- -4722
x"eb2f0",-- -5329
x"eccf0",-- -4913
x"e5190",-- -6887
x"e0330",-- -8141
x"e4c10",-- -6975
x"e5f90",-- -6663
x"e2ec0",-- -7444
x"e1000",-- -7936
x"ded80",-- -8488
x"df570",-- -8361
x"e4910",-- -7023
x"e6730",-- -6541
x"e28d0",-- -7539
x"e1e50",-- -7707
x"e5180",-- -6888
x"e9ce0",-- -5682
x"ed450",-- -4795
x"ecf00",-- -4880
x"ebf60",-- -5130
x"ed020",-- -4862
x"f20a0",-- -3574
x"f78d0",-- -2163
x"f81e0",-- -2018
x"f6d70",-- -2345
x"f6bc0",-- -2372
x"fb1a0",-- -1254
x"00c00",-- 192
x"02b20",-- 690
x"01bd0",-- 445
x"01380",-- 312
x"049b0",-- 1179
x"08c50",-- 2245
x"0aaf0",-- 2735
x"0b540",-- 2900
x"0cb80",-- 3256
x"0f810",-- 3969
x"12360",-- 4662
x"14020",-- 5122
x"158d0",-- 5517
x"18e80",-- 6376
x"172b0",-- 5931
x"152e0",-- 5422
x"19af0",-- 6575
x"1fa00",-- 8096
x"21ec0",-- 8684
x"1f8a0",-- 8074
x"1d240",-- 7460
x"206d0",-- 8301
x"22cf0",-- 8911
x"217b0",-- 8571
x"200e0",-- 8206
x"1e160",-- 7702
x"1ba80",-- 7080
x"15eb0",-- 5611
x"11540",-- 4436
x"0fb80",-- 4024
x"0eae0",-- 3758
x"09760",-- 2422
x"00030",-- 3
x"f87b0",-- -1925
x"f5d80",-- -2600
x"f71f0",-- -2273
x"f5ba0",-- -2630
x"ecd40",-- -4908
x"e7510",-- -6319
x"e5450",-- -6843
x"e6080",-- -6648
x"e7270",-- -6361
x"e4b70",-- -6985
x"e0830",-- -8061
x"e0170",-- -8169
x"e0bc0",-- -8004
x"e1090",-- -7927
x"e2fa0",-- -7430
x"e3680",-- -7320
x"e2210",-- -7647
x"e0a00",-- -8032
x"e4000",-- -7168
x"e8fa0",-- -5894
x"ea2b0",-- -5589
x"eb310",-- -5327
x"ec350",-- -5067
x"ebbb0",-- -5189
x"f1950",-- -3691
x"f7bc0",-- -2116
x"f69e0",-- -2402
x"f5dd0",-- -2595
x"f8cb0",-- -1845
x"fa940",-- -1388
x"fe820",-- -382
x"04610",-- 1121
x"02980",-- 664
x"ff830",-- -125
x"04140",-- 1044
x"08e80",-- 2280
x"0ab10",-- 2737
x"0b2e0",-- 2862
x"09f40",-- 2548
x"0b920",-- 2962
x"10c50",-- 4293
x"14fc0",-- 5372
x"141b0",-- 5147
x"13af0",-- 5039
x"18630",-- 6243
x"16ed0",-- 5869
x"178c0",-- 6028
x"1cd80",-- 7384
x"1f8f0",-- 8079
x"1fd80",-- 8152
x"1e5f0",-- 7775
x"1d190",-- 7449
x"20890",-- 8329
x"24040",-- 9220
x"239b0",-- 9115
x"1f0a0",-- 7946
x"19210",-- 6433
x"16520",-- 5714
x"16730",-- 5747
x"171a0",-- 5914
x"10cc0",-- 4300
x"06460",-- 1606
x"ffbc0",-- -68
x"fea20",-- -350
x"fd990",-- -615
x"f9610",-- -1695
x"f2060",-- -3578
x"e9bd0",-- -5699
x"e8a00",-- -5984
x"ea7e0",-- -5506
x"e82b0",-- -6101
x"e4370",-- -7113
x"e00b0",-- -8181
x"df160",-- -8426
x"e1770",-- -7817
x"e2f30",-- -7437
x"e0800",-- -8064
x"ddfb0",-- -8709
x"e02d0",-- -8147
x"e11b0",-- -7909
x"e2650",-- -7579
x"e5ec0",-- -6676
x"e4d80",-- -6952
x"e64b0",-- -6581
x"eb2c0",-- -5332
x"ec760",-- -5002
x"ed600",-- -4768
x"f1c50",-- -3643
x"f4820",-- -2942
x"f5590",-- -2727
x"f8170",-- -2025
x"fa030",-- -1533
x"fa840",-- -1404
x"fefa0",-- -262
x"02170",-- 535
x"00f20",-- 242
x"01510",-- 337
x"04d40",-- 1236
x"09170",-- 2327
x"099c0",-- 2460
x"09b80",-- 2488
x"0a300",-- 2608
x"0d6a0",-- 3434
x"12040",-- 4612
x"12390",-- 4665
x"13090",-- 4873
x"13d30",-- 5075
x"17d70",-- 6103
x"17490",-- 5961
x"16980",-- 5784
x"1b870",-- 7047
x"1e190",-- 7705
x"1f1e0",-- 7966
x"1f7d0",-- 8061
x"1d780",-- 7544
x"1e3e0",-- 7742
x"22310",-- 8753
x"24a60",-- 9382
x"21fa0",-- 8698
x"18c00",-- 6336
x"15a00",-- 5536
x"16a40",-- 5796
x"18070",-- 6151
x"143c0",-- 5180
x"089d0",-- 2205
x"ff270",-- -217
x"fe190",-- -487
x"ff740",-- -140
x"fc820",-- -894
x"f2d90",-- -3367
x"ea6c0",-- -5524
x"e8c60",-- -5946
x"e9680",-- -5784
x"e9600",-- -5792
x"e6820",-- -6526
x"e0000",-- -8192
x"ddc20",-- -8766
x"e0530",-- -8109
x"e2420",-- -7614
x"e12a0",-- -7894
x"dea10",-- -8543
x"de5b0",-- -8613
x"e0370",-- -8137
x"e2c40",-- -7484
x"e4650",-- -7067
x"e5430",-- -6845
x"e5790",-- -6791
x"e9220",-- -5854
x"ed6a0",-- -4758
x"ee710",-- -4495
x"ef510",-- -4271
x"f22b0",-- -3541
x"f5d00",-- -2608
x"f9700",-- -1680
x"fab70",-- -1353
x"f9a30",-- -1629
x"fc190",-- -999
x"018f0",-- 399
x"03630",-- 867
x"03380",-- 824
x"03f40",-- 1012
x"05600",-- 1376
x"08c30",-- 2243
x"0b950",-- 2965
x"0c9f0",-- 3231
x"0cca0",-- 3274
x"0da90",-- 3497
x"118a0",-- 4490
x"16390",-- 5689
x"14950",-- 5269
x"15820",-- 5506
x"189b0",-- 6299
x"17060",-- 5894
x"1a980",-- 6808
x"1e770",-- 7799
x"1f330",-- 7987
x"1f120",-- 7954
x"21050",-- 8453
x"204b0",-- 8267
x"205a0",-- 8282
x"22390",-- 8761
x"24470",-- 9287
x"1efb0",-- 7931
x"176f0",-- 5999
x"15030",-- 5379
x"15eb0",-- 5611
x"14690",-- 5225
x"0d740",-- 3444
x"04b80",-- 1208
x"fd760",-- -650
x"fb270",-- -1241
x"f9ec0",-- -1556
x"f6190",-- -2535
x"ef770",-- -4233
x"e8fd0",-- -5891
x"e5970",-- -6761
x"e5430",-- -6845
x"e5110",-- -6895
x"e3b60",-- -7242
x"dfdb0",-- -8229
x"ddb50",-- -8779
x"dd820",-- -8830
x"de870",-- -8569
x"dfb10",-- -8271
x"e0790",-- -8071
x"e0370",-- -8137
x"df770",-- -8329
x"e1220",-- -7902
x"e50e0",-- -6898
x"e7ea0",-- -6166
x"ea5d0",-- -5539
x"eb3e0",-- -5314
x"ec530",-- -5037
x"efbb0",-- -4165
x"f3930",-- -3181
x"f6c30",-- -2365
x"f9810",-- -1663
x"fa870",-- -1401
x"fa520",-- -1454
x"fd5d0",-- -675
x"023a0",-- 570
x"04340",-- 1076
x"03d80",-- 984
x"047b0",-- 1147
x"06670",-- 1639
x"09620",-- 2402
x"0c5a0",-- 3162
x"0d030",-- 3331
x"0d440",-- 3396
x"100a0",-- 4106
x"130e0",-- 4878
x"153b0",-- 5435
x"153a0",-- 5434
x"16f00",-- 5872
x"1bf00",-- 7152
x"182f0",-- 6191
x"183c0",-- 6204
x"1e590",-- 7769
x"222c0",-- 8748
x"23620",-- 9058
x"211a0",-- 8474
x"1dbf0",-- 7615
x"1f800",-- 8064
x"25320",-- 9522
x"26450",-- 9797
x"1ffa0",-- 8186
x"183c0",-- 6204
x"13a50",-- 5029
x"14040",-- 5124
x"155f0",-- 5471
x"0f970",-- 3991
x"04f70",-- 1271
x"fbe40",-- -1052
x"f8340",-- -1996
x"f7bc0",-- -2116
x"f6c10",-- -2367
x"f0cf0",-- -3889
x"e7520",-- -6318
x"e1db0",-- -7717
x"e2a00",-- -7520
x"e2b20",-- -7502
x"e4370",-- -7113
x"e0290",-- -8151
x"da6a0",-- -9622
x"d9660",-- -9882
x"dd950",-- -8811
x"dffe0",-- -8194
x"df4d0",-- -8371
x"df140",-- -8428
x"dce20",-- -8990
x"e0800",-- -8064
x"e6870",-- -6521
x"e7750",-- -6283
x"e85a0",-- -6054
x"ec210",-- -5087
x"ed680",-- -4760
x"f0260",-- -4058
x"f4990",-- -2919
x"f6d50",-- -2347
x"f8b10",-- -1871
x"fbf90",-- -1031
x"fd130",-- -749
x"fe750",-- -395
x"02d20",-- 722
x"04ef0",-- 1263
x"056a0",-- 1386
x"07030",-- 1795
x"08020",-- 2050
x"0a360",-- 2614
x"0cb90",-- 3257
x"0f950",-- 3989
x"10720",-- 4210
x"11d20",-- 4562
x"133d0",-- 4925
x"15820",-- 5506
x"183e0",-- 6206
x"1a900",-- 6800
x"1a640",-- 6756
x"17ee0",-- 6126
x"1b5f0",-- 7007
x"1f7d0",-- 8061
x"231a0",-- 8986
x"237e0",-- 9086
x"20730",-- 8307
x"1ecc0",-- 7884
x"213c0",-- 8508
x"247e0",-- 9342
x"24340",-- 9268
x"1e750",-- 7797
x"176f0",-- 5999
x"13040",-- 4868
x"13210",-- 4897
x"130b0",-- 4875
x"0d470",-- 3399
x"02550",-- 597
x"f9b70",-- -1609
x"f6230",-- -2525
x"f5ef0",-- -2577
x"f5950",-- -2667
x"ed4a0",-- -4790
x"e3020",-- -7422
x"df0c0",-- -8436
x"e1180",-- -7912
x"e3fe0",-- -7170
x"e2330",-- -7629
x"dc440",-- -9148
x"d79f0",-- -10337
x"d7e10",-- -10271
x"dd340",-- -8908
x"e0ab0",-- -8021
x"e0970",-- -8041
x"dc190",-- -9191
x"dafb0",-- -9477
x"e1650",-- -7835
x"e77a0",-- -6278
x"eb8b0",-- -5237
x"ebe20",-- -5150
x"e9d10",-- -5679
x"eb880",-- -5240
x"f1890",-- -3703
x"f8350",-- -1995
x"fb9e0",-- -1122
x"faad0",-- -1363
x"f94a0",-- -1718
x"fbc20",-- -1086
x"02a00",-- 672
x"06eb0",-- 1771
x"06300",-- 1584
x"05e50",-- 1509
x"082d0",-- 2093
x"09bf0",-- 2495
x"0b4f0",-- 2895
x"0dd00",-- 3536
x"0fa60",-- 4006
x"120a0",-- 4618
x"12c30",-- 4803
x"12930",-- 4755
x"15dd0",-- 5597
x"18700",-- 6256
x"1d960",-- 7574
x"1c770",-- 7287
x"175d0",-- 5981
x"1ab80",-- 6840
x"21350",-- 8501
x"25c60",-- 9670
x"25000",-- 9472
x"20220",-- 8226
x"1dad0",-- 7597
x"21690",-- 8553
x"25d20",-- 9682
x"25600",-- 9568
x"1dfa0",-- 7674
x"146b0",-- 5227
x"10230",-- 4131
x"12db0",-- 4827
x"12310",-- 4657
x"0a820",-- 2690
x"fea70",-- -345
x"f54c0",-- -2740
x"f2e60",-- -3354
x"f45c0",-- -2980
x"f1b50",-- -3659
x"e7f60",-- -6154
x"df610",-- -8351
x"dcc40",-- -9020
x"df0c0",-- -8436
x"e2530",-- -7597
x"de7d0",-- -8579
x"d8230",-- -10205
x"d5f40",-- -10764
x"d9c20",-- -9790
x"dddd0",-- -8739
x"de620",-- -8606
x"dc260",-- -9178
x"db450",-- -9403
x"df4a0",-- -8374
x"e4a10",-- -7007
x"e8b90",-- -5959
x"e9930",-- -5741
x"e92c0",-- -5844
x"eb240",-- -5340
x"f18d0",-- -3699
x"f6850",-- -2427
x"f7ce0",-- -2098
x"f87a0",-- -1926
x"f9cb0",-- -1589
x"fdb50",-- -587
x"03d60",-- 982
x"059a0",-- 1434
x"05170",-- 1303
x"05db0",-- 1499
x"08e60",-- 2278
x"0c660",-- 3174
x"0f090",-- 3849
x"0d9c0",-- 3484
x"0e1e0",-- 3614
x"11b90",-- 4537
x"15740",-- 5492
x"16720",-- 5746
x"18090",-- 6153
x"17830",-- 6019
x"1b080",-- 6920
x"1fc60",-- 8134
x"1b9e0",-- 7070
x"1b030",-- 6915
x"1d850",-- 7557
x"24190",-- 9241
x"26c70",-- 9927
x"24890",-- 9353
x"1e1d0",-- 7709
x"1d6a0",-- 7530
x"21cb0",-- 8651
x"26c50",-- 9925
x"23030",-- 8963
x"17b90",-- 6073
x"0ea50",-- 3749
x"0cf20",-- 3314
x"109f0",-- 4255
x"0ec00",-- 3776
x"05800",-- 1408
x"f6d90",-- -2343
x"ee960",-- -4458
x"eede0",-- -4386
x"f11d0",-- -3811
x"ed7a0",-- -4742
x"e3d80",-- -7208
x"da060",-- -9722
x"d83c0",-- -10180
x"dd730",-- -8845
x"dfa40",-- -8284
x"dc1f0",-- -9185
x"d6e90",-- -10519
x"d52d0",-- -10963
x"d8420",-- -10174
x"dd2f0",-- -8913
x"ddc00",-- -8768
x"dcfb0",-- -8965
x"df3e0",-- -8386
x"e1f40",-- -7692
x"e6100",-- -6640
x"e8850",-- -6011
x"e9e20",-- -5662
x"edb10",-- -4687
x"f2250",-- -3547
x"f45f0",-- -2977
x"f5dd0",-- -2595
x"f8300",-- -2000
x"fb740",-- -1164
x"00160",-- 22
x"049d0",-- 1181
x"05450",-- 1349
x"056f0",-- 1391
x"07a60",-- 1958
x"0b040",-- 2820
x"0f8d0",-- 3981
x"11e40",-- 4580
x"0fc40",-- 4036
x"0f350",-- 3893
x"12f20",-- 4850
x"17f60",-- 6134
x"19f00",-- 6640
x"1b050",-- 6917
x"1a320",-- 6706
x"1bc10",-- 7105
x"21cb0",-- 8651
x"1dd20",-- 7634
x"1d290",-- 7465
x"1f830",-- 8067
x"23710",-- 9073
x"26a20",-- 9890
x"24890",-- 9353
x"1ee80",-- 7912
x"1c930",-- 7315
x"20cf0",-- 8399
x"249f0",-- 9375
x"214c0",-- 8524
x"18310",-- 6193
x"0d6f0",-- 3439
x"099e0",-- 2462
x"0d6a0",-- 3434
x"0c700",-- 3184
x"04430",-- 1091
x"f6490",-- -2487
x"ebfe0",-- -5122
x"ea7b0",-- -5509
x"ecd00",-- -4912
x"eb2a0",-- -5334
x"e1c90",-- -7735
x"d83f0",-- -10177
x"d6e20",-- -10526
x"d8d30",-- -10029
x"dc670",-- -9113
x"dabf0",-- -9537
x"d6970",-- -10601
x"d4da0",-- -11046
x"d7f90",-- -10247
x"db220",-- -9438
x"db5f0",-- -9377
x"de1c0",-- -8676
x"e0560",-- -8106
x"e2f30",-- -7437
x"e7f60",-- -6154
x"e9ae0",-- -5714
x"ea280",-- -5592
x"eee40",-- -4380
x"f3e20",-- -3102
x"f7a80",-- -2136
x"f9bc0",-- -1604
x"f9ea0",-- -1558
x"fac60",-- -1338
x"ffe40",-- -28
x"06d10",-- 1745
x"08b60",-- 2230
x"07900",-- 1936
x"07d80",-- 2008
x"0b360",-- 2870
x"10550",-- 4181
x"13440",-- 4932
x"11970",-- 4503
x"0f8f0",-- 3983
x"134e0",-- 4942
x"18a90",-- 6313
x"19f30",-- 6643
x"1a660",-- 6758
x"19ba0",-- 6586
x"1c820",-- 7298
x"20950",-- 8341
x"1d1e0",-- 7454
x"1c3e0",-- 7230
x"1d640",-- 7524
x"22830",-- 8835
x"27000",-- 9984
x"24570",-- 9303
x"1e310",-- 7729
x"1b470",-- 6983
x"1dbe0",-- 7614
x"23380",-- 9016
x"226a0",-- 8810
x"18e50",-- 6373
x"0d0b0",-- 3339
x"07760",-- 1910
x"0a280",-- 2600
x"0ac30",-- 2755
x"052e0",-- 1326
x"f7bc0",-- -2116
x"eb630",-- -5277
x"e8190",-- -6119
x"e97e0",-- -5762
x"e9e50",-- -5659
x"e2e40",-- -7452
x"db070",-- -9465
x"d65a0",-- -10662
x"d66e0",-- -10642
x"d8e70",-- -10009
x"d8510",-- -10159
x"d7cd0",-- -10291
x"d6620",-- -10654
x"d7c00",-- -10304
x"d8dd0",-- -10019
x"d8ab0",-- -10069
x"dc170",-- -9193
x"e0ab0",-- -8021
x"e5590",-- -6823
x"e8460",-- -6074
x"e7ef0",-- -6161
x"e8100",-- -6128
x"ed290",-- -4823
x"f4c00",-- -2880
x"f9430",-- -1725
x"f9750",-- -1675
x"f9310",-- -1743
x"faca0",-- -1334
x"ffa60",-- -90
x"072e0",-- 1838
x"0acc0",-- 2764
x"09850",-- 2437
x"08aa0",-- 2218
x"0c720",-- 3186
x"11720",-- 4466
x"15010",-- 5377
x"14af0",-- 5295
x"14640",-- 5220
x"15d00",-- 5584
x"19df0",-- 6623
x"1d7d0",-- 7549
x"1e8c0",-- 7820
x"1e340",-- 7732
x"23780",-- 9080
x"23a80",-- 9128
x"1f3a0",-- 7994
x"20140",-- 8212
x"21530",-- 8531
x"27a50",-- 10149
x"2a860",-- 10886
x"25cd0",-- 9677
x"1e1d0",-- 7709
x"1bf00",-- 7152
x"1f620",-- 8034
x"22f60",-- 8950
x"1f580",-- 8024
x"15e60",-- 5606
x"093d0",-- 2365
x"042b0",-- 1067
x"066c0",-- 1644
x"05170",-- 1303
x"fdf30",-- -525
x"f1f70",-- -3593
x"e7e00",-- -6176
x"e2a30",-- -7517
x"e3ab0",-- -7253
x"e1b00",-- -7760
x"dd070",-- -8953
x"d7ae0",-- -10322
x"d5180",-- -10984
x"d3660",-- -11418
x"d2fd0",-- -11523
x"d3ef0",-- -11281
x"d4c10",-- -11071
x"d7a40",-- -10332
x"d9960",-- -9834
x"d9190",-- -9959
x"d7910",-- -10351
x"db960",-- -9322
x"e2350",-- -7627
x"e8e10",-- -5919
x"ec490",-- -5047
x"eb2a0",-- -5334
x"ea8a0",-- -5494
x"ef240",-- -4316
x"f6dc0",-- -2340
x"fce40",-- -796
x"fe4d0",-- -435
x"fe5d0",-- -419
x"febe0",-- -322
x"01e70",-- 487
x"08430",-- 2115
x"0c5f0",-- 3167
x"0d060",-- 3334
x"0de70",-- 3559
x"0f800",-- 3968
x"11800",-- 4480
x"13a60",-- 5030
x"15640",-- 5476
x"17780",-- 6008
x"1b800",-- 7040
x"1c910",-- 7313
x"1d8d0",-- 7565
x"1cbd0",-- 7357
x"21d20",-- 8658
x"261d0",-- 9757
x"20c00",-- 8384
x"21580",-- 8536
x"204d0",-- 8269
x"254b0",-- 9547
x"280c0",-- 10252
x"27ad0",-- 10157
x"1e910",-- 7825
x"18690",-- 6249
x"1d2b0",-- 7467
x"20b60",-- 8374
x"23080",-- 8968
x"198a0",-- 6538
x"09420",-- 2370
x"00990",-- 153
x"02640",-- 612
x"05dd0",-- 1501
x"00a80",-- 168
x"f4b40",-- -2892
x"e6920",-- -6510
x"de230",-- -8669
x"e2190",-- -7655
x"e3600",-- -7328
x"dfb50",-- -8267
x"da4e0",-- -9650
x"d4a60",-- -11098
x"d2ec0",-- -11540
x"d4d20",-- -11054
x"d6150",-- -10731
x"d7220",-- -10462
x"da5b0",-- -9637
x"decb0",-- -8501
x"dd000",-- -8960
x"db930",-- -9325
x"dc300",-- -9168
x"e1130",-- -7917
x"eb4a0",-- -5302
x"f2460",-- -3514
x"f1180",-- -3816
x"ec800",-- -4992
x"ee170",-- -4585
x"f4570",-- -2985
x"fddb0",-- -549
x"03f80",-- 1016
x"019f0",-- 415
x"fd590",-- -679
x"ffa80",-- -88
x"05b20",-- 1458
x"0b4e0",-- 2894
x"0ddb0",-- 3547
x"0d5e0",-- 3422
x"0cca0",-- 3274
x"0e3e0",-- 3646
x"11100",-- 4368
x"11720",-- 4466
x"13650",-- 4965
x"17330",-- 5939
x"18c20",-- 6338
x"19d20",-- 6610
x"1b030",-- 6915
x"1b350",-- 6965
x"20a10",-- 8353
x"20520",-- 8274
x"1fd80",-- 8152
x"1f710",-- 8049
x"1feb0",-- 8171
x"24db0",-- 9435
x"250f0",-- 9487
x"23960",-- 9110
x"1fff0",-- 8191
x"1e5c0",-- 7772
x"1e2d0",-- 7725
x"1ebb0",-- 7867
x"1b730",-- 7027
x"14a50",-- 5285
x"0b680",-- 2920
x"076a0",-- 1898
x"05400",-- 1344
x"01b20",-- 434
x"fc160",-- -1002
x"f1e50",-- -3611
x"ea960",-- -5482
x"e6940",-- -6508
x"e4490",-- -7095
x"e28a0",-- -7542
x"dd3c0",-- -8900
x"dad00",-- -9520
x"d7700",-- -10384
x"d73b0",-- -10437
x"d7890",-- -10359
x"d5fc0",-- -10756
x"d79a0",-- -10342
x"d8e70",-- -10009
x"dc370",-- -9161
x"dc2e0",-- -9170
x"dcfa0",-- -8966
x"de880",-- -8568
x"e2ab0",-- -7509
x"e9130",-- -5869
x"ed290",-- -4823
x"ed2a0",-- -4822
x"ee240",-- -4572
x"f0d50",-- -3883
x"f5250",-- -2779
x"fafd0",-- -1283
x"fe700",-- -400
x"ff540",-- -172
x"ffef0",-- -17
x"03810",-- 897
x"06e30",-- 1763
x"095b0",-- 2395
x"0b580",-- 2904
x"0cc30",-- 3267
x"0edb0",-- 3803
x"10e00",-- 4320
x"12590",-- 4697
x"12730",-- 4723
x"13620",-- 4962
x"16900",-- 5776
x"17dc0",-- 6108
x"1b240",-- 6948
x"1bb70",-- 7095
x"1cd90",-- 7385
x"210d0",-- 8461
x"1d760",-- 7542
x"1dff0",-- 7679
x"1f100",-- 7952
x"215d0",-- 8541
x"257e0",-- 9598
x"24a70",-- 9383
x"204b0",-- 8267
x"1dbe0",-- 7614
x"1bfa0",-- 7162
x"1db90",-- 7609
x"1e5a0",-- 7770
x"19e20",-- 6626
x"13420",-- 4930
x"09720",-- 2418
x"06500",-- 1616
x"03790",-- 889
x"fff10",-- -15
x"fb990",-- -1127
x"f2b60",-- -3402
x"ebc00",-- -5184
x"e6c90",-- -6455
x"e2e70",-- -7449
x"e06a0",-- -8086
x"de500",-- -8624
x"dcc60",-- -9018
x"da800",-- -9600
x"d8e90",-- -10007
x"d6600",-- -10656
x"d4f50",-- -11019
x"d7f40",-- -10252
x"db180",-- -9448
x"dd370",-- -8905
x"de080",-- -8696
x"dd640",-- -8860
x"deba0",-- -8518
x"e2dd0",-- -7459
x"e92c0",-- -5844
x"ec6f0",-- -5009
x"edfe0",-- -4610
x"f0b40",-- -3916
x"f2a50",-- -3419
x"f68c0",-- -2420
x"fa700",-- -1424
x"fbf90",-- -1031
x"feb90",-- -327
x"028a0",-- 650
x"06760",-- 1654
x"06b40",-- 1716
x"07c90",-- 1993
x"09b80",-- 2488
x"0c190",-- 3097
x"0e700",-- 3696
x"11ad0",-- 4525
x"117b0",-- 4475
x"0f860",-- 3974
x"116d0",-- 4461
x"12e60",-- 4838
x"184d0",-- 6221
x"18870",-- 6279
x"19bf0",-- 6591
x"1b0b0",-- 6923
x"1e450",-- 7749
x"1c6d0",-- 7277
x"1ab80",-- 6840
x"1d120",-- 7442
x"1db40",-- 7604
x"24600",-- 9312
x"250d0",-- 9485
x"21210",-- 8481
x"1c2f0",-- 7215
x"19d50",-- 6613
x"1c1d0",-- 7197
x"1d0a0",-- 7434
x"1c0f0",-- 7183
x"16540",-- 5716
x"0c430",-- 3139
x"07a60",-- 1958
x"04f90",-- 1273
x"017c0",-- 380
x"fdd10",-- -559
x"f6940",-- -2412
x"f08c0",-- -3956
x"eb790",-- -5255
x"e79d0",-- -6243
x"e4420",-- -7102
x"dfb10",-- -8271
x"df310",-- -8399
x"de050",-- -8699
x"dd370",-- -8905
x"dbca0",-- -9270
x"d8300",-- -10192
x"d8060",-- -10234
x"d9a40",-- -9820
x"de190",-- -8679
x"df360",-- -8394
x"e0230",-- -8157
x"e1090",-- -7927
x"e2a00",-- -7520
x"e6c30",-- -6461
x"eafa0",-- -5382
x"ed2a0",-- -4822
x"efc00",-- -4160
x"f3290",-- -3287
x"f5d50",-- -2603
x"f8940",-- -1900
x"fb180",-- -1256
x"fd920",-- -622
x"ff510",-- -175
x"034c0",-- 844
x"06020",-- 1538
x"071c0",-- 1820
x"076a0",-- 1898
x"09ab0",-- 2475
x"0a4a0",-- 2634
x"0e4f0",-- 3663
x"0ffa0",-- 4090
x"0d1f0",-- 3359
x"0f030",-- 3843
x"100a0",-- 4106
x"13220",-- 4898
x"13940",-- 5012
x"14660",-- 5222
x"16250",-- 5669
x"17e70",-- 6119
x"1d2b0",-- 7467
x"1c230",-- 7203
x"1a310",-- 6705
x"19670",-- 6503
x"1bd30",-- 7123
x"1fbc0",-- 8124
x"21e20",-- 8674
x"20500",-- 8272
x"1bd30",-- 7123
x"1b370",-- 6967
x"1a5a0",-- 6746
x"1a930",-- 6803
x"18430",-- 6211
x"148e0",-- 5262
x"0e930",-- 3731
x"0acc0",-- 2764
x"082d0",-- 2093
x"02710",-- 625
x"fdd80",-- -552
x"f6ad0",-- -2387
x"f4190",-- -3047
x"f0080",-- -4088
x"ed040",-- -4860
x"e8260",-- -6106
x"e22e0",-- -7634
x"e14d0",-- -7859
x"e0330",-- -8141
x"e0940",-- -8044
x"deff0",-- -8449
x"dc880",-- -9080
x"daff0",-- -9473
x"dd040",-- -8956
x"debe0",-- -8514
x"e0550",-- -8107
x"e1480",-- -7864
x"e2030",-- -7677
x"e4c10",-- -6975
x"e7fc0",-- -6148
x"eb830",-- -5245
x"ec8e0",-- -4978
x"eee30",-- -4381
x"f23f0",-- -3521
x"f5ca0",-- -2614
x"f8750",-- -1931
x"fa2f0",-- -1489
x"fc2a0",-- -982
x"fdf90",-- -519
x"01130",-- 275
x"03970",-- 919
x"03b80",-- 952
x"065a0",-- 1626
x"07cc0",-- 1996
x"06410",-- 1601
x"0c460",-- 3142
x"0a200",-- 2592
x"08fe0",-- 2302
x"0a9b0",-- 2715
x"0e190",-- 3609
x"0ea90",-- 3753
x"0ec80",-- 3784
x"14200",-- 5152
x"0f100",-- 3856
x"15350",-- 5429
x"156c0",-- 5484
x"19440",-- 6468
x"19d80",-- 6616
x"18110",-- 6161
x"19f30",-- 6643
x"19230",-- 6435
x"1e7f0",-- 7807
x"1ecc0",-- 7884
x"1db50",-- 7605
x"1a140",-- 6676
x"1b970",-- 7063
x"19080",-- 6408
x"199b0",-- 6555
x"16ca0",-- 5834
x"130d0",-- 4877
x"0f350",-- 3893
x"0b210",-- 2849
x"09c70",-- 2503
x"027d0",-- 637
x"ff7c0",-- -132
x"f9b20",-- -1614
x"f6660",-- -2458
x"f2c00",-- -3392
x"f0030",-- -4093
x"eb070",-- -5369
x"e7270",-- -6361
x"e6690",-- -6551
x"e4c10",-- -6975
x"e47d0",-- -7043
x"e1880",-- -7800
x"e11b0",-- -7909
x"ded20",-- -8494
x"e1a90",-- -7767
x"e2460",-- -7610
x"e2320",-- -7630
x"e2fb0",-- -7429
x"e3970",-- -7273
x"e7750",-- -6283
x"e97f0",-- -5761
x"eccf0",-- -4913
x"edb00",-- -4688
x"ee7d0",-- -4483
x"f1920",-- -3694
x"f4550",-- -2987
x"f7390",-- -2247
x"f99e0",-- -1634
x"fb5b0",-- -1189
x"fb940",-- -1132
x"fd470",-- -697
x"02940",-- 660
x"ff850",-- -123
x"025a0",-- 602
x"05600",-- 1376
x"04030",-- 1027
x"06f90",-- 1785
x"07030",-- 1795
x"06930",-- 1683
x"04230",-- 1059
x"0b9e0",-- 2974
x"0b3d0",-- 2877
x"090b0",-- 2315
x"0d860",-- 3462
x"0c680",-- 3176
x"0f1f0",-- 3871
x"124d0",-- 4685
x"11800",-- 4480
x"14d60",-- 5334
x"17cb0",-- 6091
x"13080",-- 4872
x"18720",-- 6258
x"17c90",-- 6089
x"17940",-- 6036
x"1c4f0",-- 7247
x"1a0e0",-- 6670
x"19d00",-- 6608
x"19640",-- 6500
x"18430",-- 6211
x"167a0",-- 5754
x"15790",-- 5497
x"12d90",-- 4825
x"114f0",-- 4431
x"0cd10",-- 3281
x"09920",-- 2450
x"070d0",-- 1805
x"01d60",-- 470
x"ffa40",-- -92
x"fa8a0",-- -1398
x"f7db0",-- -2085
x"f4dc0",-- -2852
x"f2390",-- -3527
x"eff10",-- -4111
x"ebac0",-- -5204
x"ea490",-- -5559
x"e8380",-- -6088
x"e7ef0",-- -6161
x"e62b0",-- -6613
x"e62b0",-- -6613
x"e5570",-- -6825
x"e5330",-- -6861
x"e6a10",-- -6495
x"e6ab0",-- -6485
x"e6fc0",-- -6404
x"e8af0",-- -5969
x"ea5b0",-- -5541
x"eb920",-- -5230
x"ee470",-- -4537
x"efcf0",-- -4145
x"f1700",-- -3728
x"f0260",-- -4058
x"f47d0",-- -2947
x"f4760",-- -2954
x"f6580",-- -2472
x"f9f10",-- -1551
x"f8e80",-- -1816
x"fb920",-- -1134
x"fb710",-- -1167
x"fecb0",-- -309
x"00490",-- 73
x"fce90",-- -791
x"02350",-- 565
x"057b0",-- 1403
x"ff710",-- -143
x"071f0",-- 1823
x"049d0",-- 1181
x"051f0",-- 1311
x"08580",-- 2136
x"08720",-- 2162
x"0b490",-- 2889
x"0aa40",-- 2724
x"0ea90",-- 3753
x"0db70",-- 3511
x"10bb0",-- 4283
x"11fa0",-- 4602
x"13800",-- 4992
x"12fa0",-- 4858
x"16ca0",-- 5834
x"15290",-- 5417
x"15710",-- 5489
x"15b90",-- 5561
x"13f10",-- 5105
x"19ec0",-- 6636
x"14950",-- 5269
x"17100",-- 5904
x"14ca0",-- 5322
x"13210",-- 4897
x"13b00",-- 5040
x"0f440",-- 3908
x"0f740",-- 3956
x"0b260",-- 2854
x"09f90",-- 2553
x"06140",-- 1556
x"05ae0",-- 1454
x"00c80",-- 200
x"fe5c0",-- -420
x"fb390",-- -1223
x"f80f0",-- -2033
x"f6990",-- -2407
x"f35b0",-- -3237
x"f2d90",-- -3367
x"eeaf0",-- -4433
x"ee850",-- -4475
x"ebc00",-- -5184
x"ec940",-- -4972
x"eaf80",-- -5384
x"e9860",-- -5754
x"eb0e0",-- -5362
x"e9bd0",-- -5699
x"eb930",-- -5229
x"e9ea0",-- -5654
x"eb970",-- -5225
x"eb980",-- -5224
x"ee2d0",-- -4563
x"ed5b0",-- -4773
x"f1c40",-- -3644
x"eee80",-- -4376
x"f0b70",-- -3913
x"f6d50",-- -2347
x"edc70",-- -4665
x"f8520",-- -1966
x"f5ba0",-- -2630
x"f6490",-- -2487
x"f8000",-- -2048
x"fa840",-- -1404
x"fa530",-- -1453
x"fab60",-- -1354
x"ff400",-- -192
x"f8b70",-- -1865
x"04b80",-- 1208
x"00020",-- 2
x"ffce0",-- -50
x"058d0",-- 1421
x"01d60",-- 470
x"04f20",-- 1266
x"08930",-- 2195
x"07a90",-- 1961
x"0ac80",-- 2760
x"094e0",-- 2382
x"0a680",-- 2664
x"0c7d0",-- 3197
x"0be20",-- 3042
x"11760",-- 4470
x"0e4f0",-- 3663
x"11670",-- 4455
x"0fa10",-- 4001
x"12fa0",-- 4858
x"13820",-- 4994
x"0fc10",-- 4033
x"13180",-- 4888
x"11f80",-- 4600
x"12b60",-- 4790
x"10ef0",-- 4335
x"142c0",-- 5164
x"0f810",-- 3969
x"11030",-- 4355
x"10c00",-- 4288
x"0cd90",-- 3289
x"0dc70",-- 3527
x"0aaa0",-- 2730
x"0af50",-- 2805
x"083c0",-- 2108
x"08300",-- 2096
x"03990",-- 921
x"01c90",-- 457
x"fd470",-- -697
x"fc4d0",-- -947
x"fb810",-- -1151
x"f98a0",-- -1654
x"f8700",-- -1936
x"f4160",-- -3050
x"f4050",-- -3067
x"efed0",-- -4115
x"f2280",-- -3544
x"ef1b0",-- -4325
x"f0370",-- -4041
x"ee780",-- -4488
x"ef060",-- -4346
x"ee2e0",-- -4562
x"ed750",-- -4747
x"eeed0",-- -4371
x"eb160",-- -5354
x"f0bb0",-- -3909
x"ed0e0",-- -4850
x"f34f0",-- -3249
x"ec690",-- -5015
x"f3f10",-- -3087
x"eefc0",-- -4356
x"f1d40",-- -3628
x"f5880",-- -2680
x"f0f50",-- -3851
x"fa760",-- -1418
x"f1830",-- -3709
x"fa390",-- -1479
x"f6f80",-- -2312
x"fb0b0",-- -1269
x"fa050",-- -1531
x"fc6b0",-- -917
x"fe1b0",-- -485
x"ff510",-- -175
x"008e0",-- 142
x"01db0",-- 475
x"015e0",-- 350
x"02c00",-- 704
x"05950",-- 1429
x"02aa0",-- 682
x"0a1b0",-- 2587
x"05da0",-- 1498
x"071a0",-- 1818
x"0b800",-- 2944
x"064b0",-- 1611
x"0a7d0",-- 2685
x"0c270",-- 3111
x"08e80",-- 2280
x"0f490",-- 3913
x"0cc70",-- 3271
x"0c250",-- 3109
x"109f0",-- 4255
x"0b080",-- 2824
x"12690",-- 4713
x"0e4f0",-- 3663
x"0f260",-- 3878
x"11920",-- 4498
x"0c690",-- 3177
x"11a80",-- 4520
x"0fc40",-- 4036
x"11400",-- 4416
x"0d990",-- 3481
x"0f450",-- 3909
x"0bec0",-- 3052
x"0cc50",-- 3269
x"0a9b0",-- 2715
x"0a750",-- 2677
x"08960",-- 2198
x"04260",-- 1062
x"06050",-- 1541
x"00af0",-- 175
x"01940",-- 404
x"fda10",-- -607
x"fd380",-- -712
x"f9970",-- -1641
x"f99c0",-- -1636
x"f7a40",-- -2140
x"f5070",-- -2809
x"f5430",-- -2749
x"f23c0",-- -3524
x"f30b0",-- -3317
x"f1160",-- -3818
x"f2e10",-- -3359
x"ee930",-- -4461
x"f2aa0",-- -3414
x"eeb70",-- -4425
x"ef9f0",-- -4193
x"f0990",-- -3943
x"efec0",-- -4116
x"efc40",-- -4156
x"f17e0",-- -3714
x"f3970",-- -3177
x"ef1f0",-- -4321
x"f7cb0",-- -2101
x"eea70",-- -4441
x"f74d0",-- -2227
x"f5660",-- -2714
x"f1b80",-- -3656
x"fc300",-- -976
x"f67f0",-- -2433
x"f8a20",-- -1886
x"f8570",-- -1961
x"ff590",-- -167
x"f8670",-- -1945
x"fd6c0",-- -660
x"00f00",-- 240
x"fab20",-- -1358
x"04b90",-- 1209
x"fc990",-- -871
x"05290",-- 1321
x"fdfd0",-- -515
x"05060",-- 1286
x"02460",-- 582
x"01cb0",-- 459
x"0a8b0",-- 2699
x"ffa60",-- -90
x"0b240",-- 2852
x"054a0",-- 1354
x"06ae0",-- 1710
x"0bf40",-- 3060
x"06840",-- 1668
x"0be20",-- 3042
x"0b920",-- 2962
x"0b920",-- 2962
x"0de70",-- 3559
x"0b360",-- 2870
x"0c0f0",-- 3087
x"0f220",-- 3874
x"0c3c0",-- 3132
x"0efe0",-- 3838
x"0dfa0",-- 3578
x"0d790",-- 3449
x"0ee00",-- 3808
x"0d270",-- 3367
x"0ebe0",-- 3774
x"0ca20",-- 3234
x"0e540",-- 3668
x"0a910",-- 2705
x"0c570",-- 3159
x"0b330",-- 2867
x"07a30",-- 1955
x"08000",-- 2048
x"05ad0",-- 1453
x"05760",-- 1398
x"02c00",-- 704
x"01f60",-- 502
x"fefa0",-- -262
x"ff040",-- -252
x"fb720",-- -1166
x"fb8d0",-- -1139
x"f9f40",-- -1548
x"f5560",-- -2730
x"f9130",-- -1773
x"f49d0",-- -2915
x"f3650",-- -3227
x"f59d0",-- -2659
x"f3520",-- -3246
x"f17c0",-- -3716
x"f2f70",-- -3337
x"f1740",-- -3724
x"f19f0",-- -3681
x"f3270",-- -3289
x"f0e90",-- -3863
x"f42b0",-- -3029
x"f0d50",-- -3883
x"f5330",-- -2765
x"f1c90",-- -3639
x"f45c0",-- -2980
x"f7e40",-- -2076
x"f1470",-- -3769
x"f9970",-- -1641
x"f5ce0",-- -2610
x"f5ab0",-- -2645
x"faee0",-- -1298
x"f69e0",-- -2402
x"f98d0",-- -1651
x"fb3b0",-- -1221
x"f9330",-- -1741
x"fea20",-- -350
x"fa140",-- -1516
x"ffda0",-- -38
x"fc940",-- -876
x"fda10",-- -607
x"04fe0",-- 1278
x"fbe20",-- -1054
x"03920",-- 914
x"ffd50",-- -43
x"04b80",-- 1208
x"00960",-- 150
x"03bd0",-- 957
x"05b00",-- 1456
x"03560",-- 854
x"07f60",-- 2038
x"02750",-- 629
x"0dd30",-- 3539
x"02320",-- 562
x"0af40",-- 2804
x"0a2d0",-- 2605
x"067a0",-- 1658
x"0e5a0",-- 3674
x"070d0",-- 1805
x"0cfe0",-- 3326
x"0bbf0",-- 3007
x"0c5f0",-- 3167
x"0a7c0",-- 2684
x"0f650",-- 3941
x"0a190",-- 2585
x"0c6e0",-- 3182
x"0e9f0",-- 3743
x"09060",-- 2310
x"0eae0",-- 3758
x"0c980",-- 3224
x"0b2e0",-- 2862
x"0b7c0",-- 2940
x"0a640",-- 2660
x"092b0",-- 2347
x"08cc0",-- 2252
x"063a0",-- 1594
x"05c10",-- 1473
x"05530",-- 1363
x"04440",-- 1092
x"02b10",-- 689
x"fdea0",-- -534
x"011c0",-- 284
x"fb180",-- -1256
x"fd130",-- -749
x"fc550",-- -939
x"f81e0",-- -2018
x"f9a80",-- -1624
x"f8390",-- -1991
x"f5a20",-- -2654
x"f6340",-- -2508
x"f6d40",-- -2348
x"f3750",-- -3211
x"f7570",-- -2217
x"f2eb0",-- -3349
x"f5e00",-- -2592
x"f4620",-- -2974
x"f4ff0",-- -2817
x"f3380",-- -3272
x"f4a30",-- -2909
x"f52a0",-- -2774
x"f50e0",-- -2802
x"f59d0",-- -2659
x"f51f0",-- -2785
x"f6cf0",-- -2353
x"f3bd0",-- -3139
x"f7a80",-- -2136
x"f5f10",-- -2575
x"f7400",-- -2240
x"f6f70",-- -2313
x"f7ea0",-- -2070
x"fb5b0",-- -1189
x"f5ae0",-- -2642
x"fc9d0",-- -867
x"fa490",-- -1463
x"fa990",-- -1383
x"fdbd0",-- -579
x"fc1c0",-- -996
x"ff260",-- -218
x"fbfb0",-- -1029
x"02e30",-- 739
x"fc0d0",-- -1011
x"03010",-- 769
x"008c0",-- 140
x"02d40",-- 724
x"012c0",-- 300
x"063f0",-- 1599
x"04f40",-- 1268
x"03d60",-- 982
x"06390",-- 1593
x"07540",-- 1876
x"07270",-- 1831
x"06430",-- 1603
x"0b7b0",-- 2939
x"07830",-- 1923
x"0a870",-- 2695
x"07df0",-- 2015
x"0b770",-- 2935
x"08210",-- 2081
x"09790",-- 2425
x"0d790",-- 3449
x"07760",-- 1910
x"0cea0",-- 3306
x"0b270",-- 2855
x"0a8e0",-- 2702
x"0af90",-- 2809
x"0a1c0",-- 2588
x"09fd0",-- 2557
x"07d60",-- 2006
x"0c3b0",-- 3131
x"08120",-- 2066
x"0cde0",-- 3294
x"05310",-- 1329
x"08c20",-- 2242
x"05e40",-- 1508
x"06d20",-- 1746
x"05e70",-- 1511
x"033d0",-- 829
x"04910",-- 1169
x"00640",-- 100
x"04140",-- 1044
x"fdfe0",-- -514
x"ff740",-- -140
x"fb4c0",-- -1204
x"fd2a0",-- -726
x"fab10",-- -1359
x"f9240",-- -1756
x"fcd50",-- -811
x"f6110",-- -2543
x"f95e0",-- -1698
x"f6e30",-- -2333
x"f5d00",-- -2608
x"f77c0",-- -2180
x"f4980",-- -2920
x"f6af0",-- -2385
x"f5540",-- -2732
x"f6890",-- -2423
x"f5920",-- -2670
x"f4840",-- -2940
x"f4870",-- -2937
x"f6660",-- -2458
x"f5380",-- -2760
x"f43a0",-- -3014
x"f84b0",-- -1973
x"f6910",-- -2415
x"f3130",-- -3309
x"fb990",-- -1127
x"f3a60",-- -3162
x"f8610",-- -1951
x"f7fd0",-- -2051
x"f6940",-- -2412
x"fb340",-- -1228
x"fad00",-- -1328
x"fb760",-- -1162
x"facf0",-- -1329
x"fd5d0",-- -675
x"fc8a0",-- -886
x"fc0c0",-- -1012
x"fe070",-- -505
x"02350",-- 565
x"feb90",-- -327
x"009d0",-- 157
x"03220",-- 802
x"ff0b0",-- -245
x"02640",-- 612
x"03d50",-- 981
x"03270",-- 807
x"019e0",-- 414
x"09240",-- 2340
x"06870",-- 1671
x"00f90",-- 249
x"0a070",-- 2567
x"02b40",-- 692
x"06210",-- 1569
x"096f0",-- 2415
x"03d50",-- 981
x"08f90",-- 2297
x"0a260",-- 2598
x"04f40",-- 1268
x"0a5f0",-- 2655
x"07290",-- 1833
x"063a0",-- 1594
x"09490",-- 2377
x"09cb0",-- 2507
x"09680",-- 2408
x"0bc70",-- 3015
x"08770",-- 2167
x"08140",-- 2068
x"093a0",-- 2362
x"05100",-- 1296
x"0b710",-- 2929
x"08870",-- 2183
x"08820",-- 2178
x"0b290",-- 2857
x"05330",-- 1331
x"09060",-- 2310
x"05710",-- 1393
x"03770",-- 887
x"05ee0",-- 1518
x"01f30",-- 499
x"03fe0",-- 1022
x"01db0",-- 475
x"00530",-- 83
x"fed50",-- -299
x"fe9b0",-- -357
x"fb1d0",-- -1251
x"fd590",-- -679
x"f8d70",-- -1833
x"fb9a0",-- -1126
x"fb850",-- -1147
x"f68c0",-- -2420
x"fb450",-- -1211
x"f6490",-- -2487
x"f60c0",-- -2548
x"f8eb0",-- -1813
x"f4b70",-- -2889
x"f77f0",-- -2177
x"f8b60",-- -1866
x"f5680",-- -2712
x"f5f10",-- -2575
x"f7330",-- -2253
x"f3660",-- -3226
x"f7750",-- -2187
x"f8df0",-- -1825
x"f18e0",-- -3698
x"fc1c0",-- -996
x"f6490",-- -2487
x"f71b0",-- -2277
x"f7920",-- -2158
x"f83a0",-- -1990
x"f7830",-- -2173
x"fb480",-- -1208
x"f97c0",-- -1668
x"f9330",-- -1741
x"fd310",-- -719
x"f6480",-- -2488
x"01d60",-- 470
x"f5340",-- -2764
x"008f0",-- 143
x"00020",-- 2
x"fb7b0",-- -1157
x"00f70",-- 247
x"fdfb0",-- -517
x"01600",-- 352
x"001b0",-- 27
x"02800",-- 640
x"fef00",-- -272
x"05ba0",-- 1466
x"00730",-- 115
x"02030",-- 515
x"07d10",-- 2001
x"fff60",-- -10
x"06050",-- 1541
x"04200",-- 1056
x"05630",-- 1379
x"05b70",-- 1463
x"04af0",-- 1199
x"09770",-- 2423
x"04f00",-- 1264
x"06900",-- 1680
x"07a40",-- 1956
x"05990",-- 1433
x"05cc0",-- 1484
x"09030",-- 2307
x"061b0",-- 1563
x"0b2c0",-- 2860
x"03df0",-- 991
x"09450",-- 2373
x"07830",-- 1923
x"04780",-- 1144
x"0c640",-- 3172
x"05b20",-- 1458
x"089a0",-- 2202
x"07800",-- 1920
x"05d10",-- 1489
x"05f30",-- 1523
x"097b0",-- 2427
x"05cb0",-- 1483
x"06bb0",-- 1723
x"05bc0",-- 1468
x"05440",-- 1348
x"062f0",-- 1583
x"03dd0",-- 989
x"041b0",-- 1051
x"00da0",-- 218
x"02f70",-- 759
x"fdf90",-- -519
x"02190",-- 537
x"fcf30",-- -781
x"fe0f0",-- -497
x"fde00",-- -544
x"fb150",-- -1259
x"fc7f0",-- -897
x"f8f80",-- -1800
x"fad90",-- -1319
x"f8670",-- -1945
x"f98b0",-- -1653
x"f8d50",-- -1835
x"f9790",-- -1671
x"f4cd0",-- -2867
x"f8610",-- -1951
x"f7290",-- -2263
x"f9220",-- -1758
x"f4460",-- -3002
x"fbbf0",-- -1089
x"f5b60",-- -2634
x"f5f90",-- -2567
x"fb520",-- -1198
x"f4df0",-- -2849
x"f9d50",-- -1579
x"f5ab0",-- -2645
x"fb180",-- -1256
x"f6c50",-- -2363
x"fa8f0",-- -1393
x"f8190",-- -2023
x"f91f0",-- -1761
x"fc120",-- -1006
x"f6500",-- -2480
x"ffb30",-- -77
x"f8700",-- -1936
x"ff7b0",-- -133
x"f8fd0",-- -1795
x"fc2b0",-- -981
x"fecf0",-- -305
x"fb830",-- -1149
x"009b0",-- 155
x"fc460",-- -954
x"02120",-- 530
x"fb330",-- -1229
x"03b70",-- 951
x"ff4a0",-- -182
x"00a00",-- 160
x"01c20",-- 450
x"026b0",-- 619
x"02820",-- 642
x"017c0",-- 380
x"03680",-- 872
x"01800",-- 384
x"06810",-- 1665
x"014f0",-- 335
x"07800",-- 1920
x"03400",-- 832
x"056a0",-- 1386
x"06810",-- 1665
x"024b0",-- 587
x"09ee0",-- 2542
x"026e0",-- 622
x"07590",-- 1881
x"05a90",-- 1449
x"07620",-- 1890
x"042a0",-- 1066
x"06db0",-- 1755
x"0aaa0",-- 2730
x"02a70",-- 679
x"09ea0",-- 2538
x"04530",-- 1107
x"0b130",-- 2835
x"03560",-- 854
x"09920",-- 2450
x"060c0",-- 1548
x"05f90",-- 1529
x"0a770",-- 2679
x"021c0",-- 540
x"0aea0",-- 2794
x"039a0",-- 922
x"08820",-- 2178
x"04e50",-- 1253
x"07240",-- 1828
x"052c0",-- 1324
x"017b0",-- 379
x"08aa0",-- 2218
x"fca70",-- -857
x"069a0",-- 1690
x"ff240",-- -220
x"ff630",-- -157
x"01f60",-- 502
x"fbf40",-- -1036
x"fe610",-- -415
x"faaa0",-- -1366
x"fbd10",-- -1071
x"f96a0",-- -1686
x"fe430",-- -445
x"f6980",-- -2408
x"fa580",-- -1448
x"fa8a0",-- -1398
x"f3a10",-- -3167
x"fa340",-- -1484
x"f82a0",-- -2006
x"f7830",-- -2173
x"f82d0",-- -2003
x"f8300",-- -2000
x"f49d0",-- -2915
x"fc190",-- -999
x"f3e00",-- -3104
x"f9770",-- -1673
x"fae90",-- -1303
x"f4bb0",-- -2885
x"fd790",-- -647
x"f47b0",-- -2949
x"fba90",-- -1111
x"f7a20",-- -2142
x"f8300",-- -2000
x"fcb40",-- -844
x"f83a0",-- -1990
x"fc6e0",-- -914
x"fd150",-- -747
x"f7c40",-- -2108
x"fc550",-- -939
x"feb20",-- -334
x"f7fb0",-- -2053
x"01c60",-- 454
x"fcaa0",-- -854
x"fbf60",-- -1034
x"00cd0",-- 205
x"fc210",-- -991
x"fff10",-- -15
x"009e0",-- 158
x"fd130",-- -749
x"04db0",-- 1243
x"00af0",-- 175
x"fde40",-- -540
x"08250",-- 2085
x"fd2a0",-- -726
x"03450",-- 837
x"04f90",-- 1273
x"01a90",-- 425
x"03880",-- 904
x"04dc0",-- 1244
x"04d20",-- 1234
x"055d0",-- 1373
x"02ad0",-- 685
x"058b0",-- 1419
x"07330",-- 1843
x"04960",-- 1174
x"073f0",-- 1855
x"09740",-- 2420
x"01860",-- 390
x"09d10",-- 2513
x"05bc0",-- 1468
x"04990",-- 1177
x"0acc0",-- 2764
x"05ec0",-- 1516
x"09270",-- 2343
x"04200",-- 1056
x"0b180",-- 2840
x"07860",-- 1926
x"06de0",-- 1758
x"0ba10",-- 2977
x"04910",-- 1169
x"0a200",-- 2592
x"08960",-- 2198
x"0a2a0",-- 2602
x"07a60",-- 1958
x"07470",-- 1863
x"0adb0",-- 2779
x"02f40",-- 756
x"08440",-- 2116
x"053f0",-- 1343
x"06a50",-- 1701
x"014f0",-- 335
x"02e00",-- 736
x"02ed0",-- 749
x"fcd40",-- -812
x"01f10",-- 497
x"fa2a0",-- -1494
x"fed90",-- -295
x"f9e50",-- -1563
x"fab70",-- -1353
x"fac30",-- -1341
x"f8250",-- -2011
x"f96f0",-- -1681
x"f7590",-- -2215
x"f9fb0",-- -1541
x"f5a60",-- -2650
x"f8d50",-- -1835
x"f6780",-- -2440
x"f6d70",-- -2345
x"f5470",-- -2745
x"fa7a0",-- -1414
x"f4ed0",-- -2835
x"f76b0",-- -2197
x"fad50",-- -1323
x"f4f00",-- -2832
x"fa4e0",-- -1458
x"f7060",-- -2298
x"f9310",-- -1743
x"f7430",-- -2237
x"fa140",-- -1516
x"f8520",-- -1966
x"f92f0",-- -1745
x"fc8f0",-- -881
x"f7290",-- -2263
x"fbf60",-- -1034
x"f7f80",-- -2056
x"fbc70",-- -1081
x"fd740",-- -652
x"f9380",-- -1736
x"f96b0",-- -1685
x"ff6d0",-- -147
x"fa530",-- -1453
x"fee40",-- -284
x"fc460",-- -954
x"fbbd0",-- -1091
x"03040",-- 772
x"fa9d0",-- -1379
x"02f20",-- 754
x"fa640",-- -1436
x"08db0",-- 2267
x"fa210",-- -1503
x"023e0",-- 574
x"02f50",-- 757
x"fd4c0",-- -692
x"06f90",-- 1785
x"019a0",-- 410
x"05fe0",-- 1534
x"ffad0",-- -83
x"08b30",-- 2227
x"fee80",-- -280
x"056d0",-- 1389
x"07a30",-- 1955
x"059c0",-- 1436
x"051d0",-- 1309
x"06580",-- 1624
x"092e0",-- 2350
x"03710",-- 881
x"058d0",-- 1421
x"09900",-- 2448
x"07f90",-- 2041
x"06980",-- 1688
x"0b8b0",-- 2955
x"060f0",-- 1551
x"09450",-- 2373
x"0a1c0",-- 2588
x"07a80",-- 1960
x"0df10",-- 3569
x"06530",-- 1619
x"0b9e0",-- 2974
x"07f10",-- 2033
x"0adb0",-- 2779
x"0d5d0",-- 3421
x"06170",-- 1559
x"0c660",-- 3174
x"07490",-- 1865
x"09030",-- 2307
x"09030",-- 2307
x"09ea0",-- 2538
x"023c0",-- 572
x"06690",-- 1641
x"03880",-- 904
x"01100",-- 272
x"04e30",-- 1251
x"fdb80",-- -584
x"00710",-- 113
x"fade0",-- -1314
x"f9e40",-- -1564
x"faed0",-- -1299
x"f9a80",-- -1624
x"f7400",-- -2240
x"f7810",-- -2175
x"f72f0",-- -2257
x"f7160",-- -2282
x"f4710",-- -2959
x"f56d0",-- -2707
x"f56d0",-- -2707
x"f52a0",-- -2774
x"f7f40",-- -2060
x"f42b0",-- -3029
x"f7400",-- -2240
x"f4ca0",-- -2870
x"f55c0",-- -2724
x"f7d10",-- -2095
x"f8890",-- -1911
x"f6530",-- -2477
x"f7ce0",-- -2098
x"f97c0",-- -1668
x"f6c10",-- -2367
x"faf70",-- -1289
x"f7750",-- -2187
x"f7400",-- -2240
x"fc070",-- -1017
x"fa870",-- -1401
x"f4230",-- -3037
x"015b0",-- 347
x"f8c30",-- -1853
x"f4370",-- -3017
x"fd900",-- -624
x"fbe00",-- -1056
x"f8ac0",-- -1876
x"fdef0",-- -529
x"ff860",-- -122
x"f9610",-- -1695
x"fc5c0",-- -932
x"ff4f0",-- -177
x"fde70",-- -537
x"fd020",-- -766
x"03210",-- 801
x"fd5b0",-- -677
x"05310",-- 1329
x"fb130",-- -1261
x"06db0",-- 1755
x"00070",-- 7
x"fe660",-- -410
x"0dc40",-- 3524
x"fb010",-- -1279
x"07940",-- 1940
x"049b0",-- 1179
x"fd5d0",-- -675
x"09490",-- 2377
x"06cd0",-- 1741
x"fe990",-- -359
x"09ea0",-- 2538
x"05b30",-- 1459
x"02490",-- 585
x"096c0",-- 2412
x"086b0",-- 2155
x"05db0",-- 1499
x"08ed0",-- 2285
x"06ae0",-- 1710
x"0c180",-- 3096
x"03d50",-- 981
x"0f5e0",-- 3934
x"0ac80",-- 2760
x"04780",-- 1144
x"17830",-- 6019
x"03e40",-- 996
x"0c4d0",-- 3149
x"11f00",-- 4592
x"08fc0",-- 2300
x"0cfc0",-- 3324
x"12a20",-- 4770
x"0aea0",-- 2794
x"0ba30",-- 2979
x"0f1c0",-- 3868
x"07e50",-- 2021
x"0dec0",-- 3564
x"06890",-- 1673
x"07950",-- 1941
x"061e0",-- 1566
x"ffd50",-- -43
x"04a00",-- 1184
x"fdc90",-- -567
x"fe080",-- -504
x"fb480",-- -1208
x"f6f00",-- -2320
x"f8570",-- -1961
x"f7830",-- -2173
x"f40f0",-- -3057
x"f44d0",-- -2995
x"f2760",-- -3466
x"f2230",-- -3549
x"f2cb0",-- -3381
x"f01f0",-- -4065
x"f5d10",-- -2607
x"f0d40",-- -3884
x"f36f0",-- -3217
x"f3720",-- -3214
x"f2870",-- -3449
x"f6670",-- -2457
x"f34d0",-- -3251
x"f8260",-- -2010
x"f5b10",-- -2639
x"f70b0",-- -2293
x"f9650",-- -1691
x"f7200",-- -2272
x"f8610",-- -1951
x"f95c0",-- -1700
x"f72a0",-- -2262
x"fc910",-- -879
x"f7f30",-- -2061
x"fcd90",-- -807
x"fa3f0",-- -1473
x"f3450",-- -3259
x"ffb20",-- -78
x"f8d90",-- -1831
x"f91d0",-- -1763
x"fbba0",-- -1094
x"fb430",-- -1213
x"fb810",-- -1151
x"f8e80",-- -1816
x"fad40",-- -1324
x"ffa60",-- -90
x"f72f0",-- -2257
x"feff0",-- -257
x"00480",-- 72
x"fbe90",-- -1047
x"03130",-- 787
x"fc6e0",-- -914
x"fcac0",-- -852
x"05830",-- 1411
x"fc570",-- -937
x"00500",-- 80
x"05e20",-- 1506
x"03360",-- 822
x"ff380",-- -200
x"09ee0",-- 2542
x"fc980",-- -872
x"06900",-- 1680
x"095e0",-- 2398
x"fd7e0",-- -642
x"13310",-- 4913
x"ffd10",-- -47
x"09f80",-- 2552
x"08120",-- 2066
x"02cc0",-- 716
x"0f3b0",-- 3899
x"05760",-- 1398
x"0dff0",-- 3583
x"0b3b0",-- 2875
x"09010",-- 2305
x"13510",-- 4945
x"07620",-- 1890
x"0cfe0",-- 3326
x"11fb0",-- 4603
x"119e0",-- 4510
x"0ed70",-- 3799
x"0d790",-- 3449
x"10220",-- 4130
x"0e980",-- 3736
x"118f0",-- 4495
x"0f350",-- 3893
x"12b80",-- 4792
x"10e60",-- 4326
x"08250",-- 2085
x"11cb0",-- 4555
x"08320",-- 2098
x"09270",-- 2343
x"08b10",-- 2225
x"ffcc0",-- -52
x"06fe0",-- 1790
x"fe160",-- -490
x"fc960",-- -874
x"f9c60",-- -1594
x"f5da0",-- -2598
x"f51b0",-- -2789
x"f39d0",-- -3171
x"f3970",-- -3177
x"f1c00",-- -3648
x"eda70",-- -4697
x"ee3a0",-- -4550
x"eef00",-- -4368
x"ed3e0",-- -4802
x"efe80",-- -4120
x"ef630",-- -4253
x"f0980",-- -3944
x"f0010",-- -4095
x"f1790",-- -3719
x"f2e90",-- -3351
x"f3070",-- -3321
x"f3b00",-- -3152
x"f63c0",-- -2500
x"f7ec0",-- -2068
x"f73e0",-- -2242
x"f8f20",-- -1806
x"f8cf0",-- -1841
x"f89e0",-- -1890
x"fb360",-- -1226
x"faa30",-- -1373
x"fa0c0",-- -1524
x"fc3c0",-- -964
x"f9fe0",-- -1538
x"f84b0",-- -1973
x"fdda0",-- -550
x"fc0a0",-- -1014
x"fa070",-- -1529
x"faff0",-- -1281
x"f82d0",-- -2003
x"fd440",-- -700
x"f8d90",-- -1831
x"faeb0",-- -1301
x"fab10",-- -1359
x"f71d0",-- -2275
x"fc6e0",-- -914
x"faad0",-- -1363
x"fd150",-- -747
x"fd0b0",-- -757
x"fc980",-- -872
x"00340",-- 52
x"fb310",-- -1231
x"01810",-- 385
x"024e0",-- 590
x"008f0",-- 143
x"02140",-- 532
x"02bb0",-- 699
x"04e00",-- 1248
x"00af0",-- 175
x"081b0",-- 2075
x"07dd0",-- 2013
x"035d0",-- 861
x"0da40",-- 3492
x"0acf0",-- 2767
x"01090",-- 265
x"102a0",-- 4138
x"08a20",-- 2210
x"0bf10",-- 3057
x"11300",-- 4400
x"09ef0",-- 2543
x"11720",-- 4466
x"0a900",-- 2704
x"12110",-- 4625
x"14020",-- 5122
x"12780",-- 4728
x"15640",-- 5476
x"13f80",-- 5112
x"10b10",-- 4273
x"0e8c0",-- 3724
x"18a20",-- 6306
x"14cd0",-- 5325
x"15cb0",-- 5579
x"14c50",-- 5317
x"10780",-- 4216
x"10e00",-- 4320
x"0dc10",-- 3521
x"11400",-- 4416
x"0b510",-- 2897
x"08080",-- 2056
x"06ed0",-- 1773
x"ffec0",-- -20
x"ff400",-- -192
x"fc050",-- -1019
x"f67a0",-- -2438
x"f60d0",-- -2547
x"f2c80",-- -3384
x"ef040",-- -4348
x"efea0",-- -4118
x"ea170",-- -5609
x"eaee0",-- -5394
x"e92e0",-- -5842
x"ea230",-- -5597
x"eb970",-- -5225
x"ea490",-- -5559
x"e9220",-- -5854
x"ea5f0",-- -5537
x"ebce0",-- -5170
x"ecbe0",-- -4930
x"effc0",-- -4100
x"ef310",-- -4303
x"f1f60",-- -3594
x"f2230",-- -3549
x"f5590",-- -2727
x"f6b10",-- -2383
x"f7540",-- -2220
x"f8260",-- -2010
x"f8dc0",-- -1828
x"f9d50",-- -1579
x"fbc40",-- -1084
x"fd670",-- -665
x"fc700",-- -912
x"fccf0",-- -817
x"fd990",-- -615
x"fd6a0",-- -662
x"008e0",-- 142
x"fe760",-- -394
x"fe850",-- -379
x"fc1c0",-- -996
x"fee30",-- -285
x"fe000",-- -512
x"fba40",-- -1116
x"ff4e0",-- -178
x"fc5c0",-- -932
x"fdc40",-- -572
x"fe4b0",-- -437
x"fb0b0",-- -1269
x"fbfd0",-- -1027
x"fe3e0",-- -450
x"fd9f0",-- -609
x"fe530",-- -429
x"ff3a0",-- -198
x"fbf40",-- -1036
x"fe640",-- -412
x"ff800",-- -128
x"00c80",-- 200
x"03bc0",-- 956
x"ff940",-- -108
x"03f80",-- 1016
x"01670",-- 359
x"053f0",-- 1343
x"07c70",-- 1991
x"07fd0",-- 2045
x"08b40",-- 2228
x"098d0",-- 2445
x"0c4a0",-- 3146
x"0b8f0",-- 2959
x"0dd30",-- 3539
x"0e0e0",-- 3598
x"104f0",-- 4175
x"10e30",-- 4323
x"117e0",-- 4478
x"159b0",-- 5531
x"14540",-- 5204
x"152b0",-- 5419
x"1b190",-- 6937
x"182d0",-- 6189
x"0f9c0",-- 3996
x"148b0",-- 5259
x"18a20",-- 6306
x"18b30",-- 6323
x"19640",-- 6500
x"16aa0",-- 5802
x"12090",-- 4617
x"0e000",-- 3584
x"0f510",-- 3921
x"10fa0",-- 4346
x"10140",-- 4116
x"083a0",-- 2106
x"02c60",-- 710
x"ff470",-- -185
x"fbbf0",-- -1089
x"fa1c0",-- -1508
x"f76a0",-- -2198
x"f2f50",-- -3339
x"ef880",-- -4216
x"eb8b0",-- -5237
x"e9b80",-- -5704
x"e8880",-- -6008
x"e4e20",-- -6942
x"e5930",-- -6765
x"e88c0",-- -6004
x"e8230",-- -6109
x"e79f0",-- -6241
x"e5540",-- -6828
x"e6730",-- -6541
x"e8aa0",-- -5974
x"ebfe0",-- -5122
x"ef7a0",-- -4230
x"efe30",-- -4125
x"eea70",-- -4441
x"eea00",-- -4448
x"f3590",-- -3239
x"f65f0",-- -2465
x"f7a90",-- -2135
x"f9240",-- -1756
x"f9d00",-- -1584
x"f9e90",-- -1559
x"fac10",-- -1343
x"fc690",-- -919
x"fd3d0",-- -707
x"fe850",-- -379
x"fff90",-- -7
x"00e80",-- 232
x"febc0",-- -324
x"fbbf0",-- -1089
x"fcfc0",-- -772
x"ffe50",-- -27
x"01ec0",-- 492
x"01cc0",-- 460
x"feb60",-- -330
x"fa640",-- -1436
x"fc5f0",-- -929
x"fe4d0",-- -435
x"00c80",-- 200
x"fff40",-- -12
x"fce60",-- -794
x"fd990",-- -615
x"fda10",-- -607
x"fd010",-- -767
x"ff8a0",-- -118
x"ffcc0",-- -52
x"feb10",-- -335
x"01c70",-- 455
x"01d50",-- 469
x"001e0",-- 30
x"01150",-- 277
x"035e0",-- 862
x"04fc0",-- 1276
x"074a0",-- 1866
x"09740",-- 2420
x"06b60",-- 1718
x"08d20",-- 2258
x"0a890",-- 2697
x"0b810",-- 2945
x"0ffa0",-- 4090
x"11290",-- 4393
x"0fae0",-- 4014
x"10540",-- 4180
x"14770",-- 5239
x"17010",-- 5889
x"1aa00",-- 6816
x"1b0f0",-- 6927
x"19bf0",-- 6591
x"151f0",-- 5407
x"14090",-- 5129
x"182c0",-- 6188
x"1d6c0",-- 7532
x"1fa00",-- 8096
x"19380",-- 6456
x"16450",-- 5701
x"121d0",-- 4637
x"10230",-- 4131
x"15ba0",-- 5562
x"12730",-- 4723
x"0c730",-- 3187
x"05e90",-- 1513
x"fec10",-- -319
x"fda40",-- -604
x"fa110",-- -1519
x"f7400",-- -2240
x"f3e70",-- -3097
x"ef680",-- -4248
x"ead00",-- -5424
x"e6f10",-- -6415
x"e5f90",-- -6663
x"e3ba0",-- -7238
x"e3320",-- -7374
x"e5ca0",-- -6710
x"e66f0",-- -6545
x"e3c00",-- -7232
x"e1a10",-- -7775
x"e28c0",-- -7540
x"e5e30",-- -6685
x"e9720",-- -5774
x"ec690",-- -5015
x"ec990",-- -4967
x"eaf30",-- -5389
x"eb970",-- -5225
x"f09d0",-- -3939
x"f58b0",-- -2677
x"f6cd0",-- -2355
x"f71a0",-- -2278
x"f7f10",-- -2063
x"f7d80",-- -2088
x"f8670",-- -1945
x"fc5c0",-- -932
x"fe7f0",-- -385
x"00120",-- 18
x"fff30",-- -13
x"ff1f0",-- -225
x"ff8d0",-- -115
x"ff0e0",-- -242
x"01970",-- 407
x"03c20",-- 962
x"03bc0",-- 956
x"01e00",-- 480
x"00eb0",-- 235
x"fe0a0",-- -502
x"fe5a0",-- -422
x"02f00",-- 752
x"02f50",-- 757
x"03e40",-- 996
x"fee40",-- -284
x"fb4f0",-- -1201
x"fef50",-- -267
x"01150",-- 277
x"01310",-- 305
x"020f0",-- 527
x"fe340",-- -460
x"fb7b0",-- -1157
x"fe570",-- -425
x"00110",-- 17
x"02190",-- 537
x"02410",-- 577
x"01940",-- 404
x"00e10",-- 225
x"03630",-- 867
x"04500",-- 1104
x"06140",-- 1556
x"0a3c0",-- 2620
x"08cd0",-- 2253
x"0be50",-- 3045
x"0bea0",-- 3050
x"0cae0",-- 3246
x"11240",-- 4388
x"11f80",-- 4600
x"15fb0",-- 5627
x"180f0",-- 6159
x"165a0",-- 5722
x"1a4b0",-- 6731
x"1b0b0",-- 6923
x"15560",-- 5462
x"17100",-- 5904
x"1b2b0",-- 6955
x"1d8f0",-- 7567
x"1ea40",-- 7844
x"1af20",-- 6898
x"159b0",-- 5531
x"13be0",-- 5054
x"13270",-- 4903
x"15730",-- 5491
x"14050",-- 5125
x"0c730",-- 3187
x"02280",-- 552
x"fdf60",-- -522
x"fe460",-- -442
x"fc280",-- -984
x"f9a40",-- -1628
x"f39d0",-- -3171
x"ece60",-- -4890
x"e7cf0",-- -6193
x"e74f0",-- -6321
x"e81f0",-- -6113
x"e6690",-- -6551
x"e3db0",-- -7205
x"e42b0",-- -7125
x"e3ab0",-- -7253
x"e2010",-- -7679
x"e2af0",-- -7505
x"e43a0",-- -7110
x"e7430",-- -6333
x"e9bf0",-- -5697
x"eb390",-- -5319
x"ea5b0",-- -5541
x"ea6e0",-- -5522
x"ec440",-- -5052
x"f14f0",-- -3761
x"f6de0",-- -2338
x"f6be0",-- -2370
x"f4fa0",-- -2822
x"f4b70",-- -2889
x"f6bb0",-- -2373
x"fa870",-- -1401
x"fd440",-- -700
x"fdbd0",-- -579
x"fd3f0",-- -705
x"fced0",-- -787
x"00190",-- 25
x"01450",-- 325
x"00df0",-- 223
x"01d80",-- 472
x"021c0",-- 540
x"03360",-- 822
x"03df0",-- 991
x"02730",-- 627
x"01680",-- 360
x"00d70",-- 215
x"01f40",-- 500
x"04a50",-- 1189
x"03590",-- 857
x"ffdd0",-- -35
x"fe250",-- -475
x"fea30",-- -349
x"00a50",-- 165
x"023e0",-- 574
x"017b0",-- 379
x"fe700",-- -400
x"fd4f0",-- -689
x"fe670",-- -409
x"00140",-- 20
x"01f60",-- 502
x"00c80",-- 200
x"ffc10",-- -63
x"019a0",-- 410
x"01b00",-- 432
x"038f0",-- 911
x"05240",-- 1316
x"05db0",-- 1499
x"09150",-- 2325
x"09970",-- 2455
x"09f10",-- 2545
x"0af90",-- 2809
x"0d210",-- 3361
x"0f510",-- 3921
x"140c0",-- 5132
x"161b0",-- 5659
x"14b90",-- 5305
x"17920",-- 6034
x"1a090",-- 6665
x"16820",-- 5762
x"16950",-- 5781
x"184a0",-- 6218
x"18c20",-- 6338
x"201e0",-- 8222
x"1e6b0",-- 7787
x"17ee0",-- 6126
x"145f0",-- 5215
x"11260",-- 4390
x"143c0",-- 5180
x"16e10",-- 5857
x"13010",-- 4865
x"09260",-- 2342
x"fef30",-- -269
x"fcfc0",-- -772
x"ff560",-- -170
x"feb90",-- -327
x"f8f80",-- -1800
x"f0460",-- -4026
x"e9890",-- -5751
x"e5e50",-- -6683
x"e85d0",-- -6051
x"eacb0",-- -5429
x"e7ab0",-- -6229
x"e4580",-- -7080
x"e2420",-- -7614
x"e2320",-- -7630
x"e3740",-- -7308
x"e4670",-- -7065
x"e74d0",-- -6323
x"e9a20",-- -5726
x"e9420",-- -5822
x"e9290",-- -5847
x"e9470",-- -5817
x"eaaf0",-- -5457
x"eeed0",-- -4371
x"f4120",-- -3054
x"f6ed0",-- -2323
x"f3c50",-- -3131
x"f1d10",-- -3631
x"f4710",-- -2959
x"f8be0",-- -1858
x"fcda0",-- -806
x"fedf0",-- -289
x"fc890",-- -887
x"f8ac0",-- -1876
x"fb3e0",-- -1218
x"001c0",-- 28
x"04610",-- 1121
x"04940",-- 1172
x"01130",-- 275
x"007d0",-- 125
x"01ad0",-- 429
x"04340",-- 1076
x"06250",-- 1573
x"066c0",-- 1644
x"02200",-- 544
x"00e80",-- 232
x"042b0",-- 1067
x"03a10",-- 929
x"04940",-- 1172
x"02ad0",-- 685
x"00800",-- 128
x"016a0",-- 362
x"00e80",-- 232
x"00c50",-- 197
x"00490",-- 73
x"fd9e0",-- -610
x"fde70",-- -537
x"ffef0",-- -17
x"ff670",-- -153
x"fd4c0",-- -692
x"fd3f0",-- -705
x"fdae0",-- -594
x"febe0",-- -322
x"01b30",-- 435
x"01b30",-- 435
x"01d00",-- 464
x"02390",-- 569
x"03e70",-- 999
x"08340",-- 2100
x"09620",-- 2402
x"096c0",-- 2412
x"0c310",-- 3121
x"0d9e0",-- 3486
x"10e50",-- 4325
x"12f90",-- 4857
x"13cd0",-- 5069
x"176c0",-- 5996
x"19b40",-- 6580
x"19ff0",-- 6655
x"19580",-- 6488
x"16390",-- 5689
x"15030",-- 5379
x"1b580",-- 7000
x"20450",-- 8261
x"1f1a0",-- 7962
x"17b20",-- 6066
x"10640",-- 4196
x"117b0",-- 4475
x"13dd0",-- 5085
x"152e0",-- 5422
x"11c40",-- 4548
x"05f60",-- 1526
x"fcd90",-- -807
x"fcde0",-- -802
x"feb60",-- -330
x"fc890",-- -887
x"f7510",-- -2223
x"eeed0",-- -4371
x"e8510",-- -6063
x"e8240",-- -6108
x"e9ce0",-- -5682
x"ea030",-- -5629
x"e82b0",-- -6101
x"e5310",-- -6863
x"e38b0",-- -7285
x"e4b40",-- -6988
x"e4dc0",-- -6948
x"e5d60",-- -6698
x"e8e90",-- -5911
x"ea820",-- -5502
x"eb0c0",-- -5364
x"ea300",-- -5584
x"ea260",-- -5594
x"ec5a0",-- -5030
x"f0cf0",-- -3889
x"f5100",-- -2800
x"f5f30",-- -2573
x"f3380",-- -3272
x"f1c70",-- -3641
x"f4f70",-- -2825
x"fad50",-- -1323
x"fd1b0",-- -741
x"fd560",-- -682
x"fbda0",-- -1062
x"fa320",-- -1486
x"fbe40",-- -1052
x"ffee0",-- -18
x"042d0",-- 1069
x"04a50",-- 1189
x"02ca0",-- 714
x"00ed0",-- 237
x"00e40",-- 228
x"031d0",-- 797
x"05630",-- 1379
x"061c0",-- 1564
x"06050",-- 1541
x"02a80",-- 680
x"00a00",-- 160
x"00c80",-- 200
x"027b0",-- 635
x"052c0",-- 1324
x"03fd0",-- 1021
x"00340",-- 52
x"fce90",-- -791
x"fbc90",-- -1079
x"ff3b0",-- -197
x"01bf0",-- 447
x"018a0",-- 394
x"fe250",-- -475
x"faf80",-- -1288
x"fb6f0",-- -1169
x"fdb80",-- -584
x"014c0",-- 332
x"018f0",-- 399
x"ff9f0",-- -97
x"feaa0",-- -342
x"ff2e0",-- -210
x"01ba0",-- 442
x"05c40",-- 1476
x"084b0",-- 2123
x"08170",-- 2071
x"07b80",-- 1976
x"09670",-- 2407
x"0b940",-- 2964
x"0f810",-- 3969
x"114e0",-- 4430
x"13a80",-- 5032
x"169b0",-- 5787
x"155d0",-- 5469
x"17cd0",-- 6093
x"1ad40",-- 6868
x"17dc0",-- 6108
x"16f40",-- 5876
x"18890",-- 6281
x"1bb00",-- 7088
x"1e7f0",-- 7807
x"1b3c0",-- 6972
x"15030",-- 5379
x"11010",-- 4353
x"12dc0",-- 4828
x"16810",-- 5761
x"12ed0",-- 4845
x"0b4c0",-- 2892
x"02bc0",-- 700
x"fdf90",-- -519
x"fe960",-- -362
x"fffb0",-- -5
x"fc210",-- -991
x"f2840",-- -3452
x"ebe70",-- -5145
x"e9cf0",-- -5681
x"eaf20",-- -5390
x"ec460",-- -5050
x"ea4c0",-- -5556
x"e6ba0",-- -6470
x"e4460",-- -7098
x"e3ce0",-- -7218
x"e65a0",-- -6566
x"e7a90",-- -6231
x"e79c0",-- -6244
x"e8e10",-- -5919
x"ea8f0",-- -5489
x"eaa60",-- -5466
x"e9830",-- -5757
x"eae40",-- -5404
x"ef510",-- -4271
x"f2ad0",-- -3411
x"f43a0",-- -3014
x"f2d20",-- -3374
x"f1bd0",-- -3651
x"f3070",-- -3321
x"f79f0",-- -2145
x"fd4c0",-- -692
x"fd600",-- -672
x"f9ab0",-- -1621
x"f88c0",-- -1908
x"fc2d0",-- -979
x"00f90",-- 249
x"03510",-- 849
x"01180",-- 280
x"ffcc0",-- -52
x"01620",-- 354
x"04850",-- 1157
x"062d0",-- 1581
x"04bb0",-- 1211
x"03080",-- 776
x"03d60",-- 982
x"05ef0",-- 1519
x"059c0",-- 1436
x"038f0",-- 911
x"00640",-- 100
x"ff4e0",-- -178
x"045c0",-- 1116
x"05860",-- 1414
x"00cf0",-- 207
x"fcbe0",-- -834
x"fa750",-- -1419
x"fe2d0",-- -467
x"02960",-- 662
x"00760",-- 118
x"fc550",-- -939
x"f8d50",-- -1835
x"f98b0",-- -1653
x"feb90",-- -327
x"01fd0",-- 509
x"ff600",-- -160
x"fb710",-- -1167
x"fc280",-- -984
x"ff620",-- -158
x"03270",-- 807
x"04f20",-- 1266
x"04280",-- 1064
x"040d0",-- 1037
x"06610",-- 1633
x"0a840",-- 2692
x"0d740",-- 3444
x"0d990",-- 3481
x"0e9b0",-- 3739
x"10b80",-- 4280
x"149d0",-- 5277
x"16b40",-- 5812
x"17dd0",-- 6109
x"19370",-- 6455
x"19470",-- 6471
x"1adc0",-- 6876
x"18410",-- 6209
x"17c60",-- 6086
x"1e7d0",-- 7805
x"1fe70",-- 8167
x"1c360",-- 7222
x"15540",-- 5460
x"11450",-- 4421
x"15d20",-- 5586
x"16050",-- 5637
x"10fa0",-- 4346
x"0c220",-- 3106
x"03b30",-- 947
x"fcaa0",-- -854
x"fd3d0",-- -707
x"014e0",-- 334
x"fb650",-- -1179
x"efd40",-- -4140
x"ebf70",-- -5129
x"ea300",-- -5584
x"ea3f0",-- -5569
x"eb130",-- -5357
x"ea490",-- -5559
x"e7660",-- -6298
x"e2850",-- -7547
x"e25b0",-- -7589
x"e7130",-- -6381
x"e86c0",-- -6036
x"e78e0",-- -6258
x"e88d0",-- -6003
x"ea960",-- -5482
x"e8ab0",-- -5973
x"e7740",-- -6284
x"ed4a0",-- -4790
x"f1890",-- -3703
x"f2080",-- -3576
x"f18b0",-- -3701
x"f1c50",-- -3643
x"f2370",-- -3529
x"f3700",-- -3216
x"f9d50",-- -1579
x"fe5a0",-- -422
x"fa9e0",-- -1378
x"f83a0",-- -1990
x"faa30",-- -1373
x"fdb20",-- -590
x"01220",-- 290
x"042a0",-- 1066
x"046b0",-- 1131
x"00530",-- 83
x"fd240",-- -732
x"03150",-- 789
x"0a5f0",-- 2655
x"0a7d0",-- 2685
x"056a0",-- 1386
x"01d30",-- 467
x"01090",-- 265
x"02050",-- 517
x"09260",-- 2342
x"0a6d0",-- 2669
x"03290",-- 809
x"fbef0",-- -1041
x"fa9d0",-- -1379
x"01220",-- 290
x"04200",-- 1056
x"021c0",-- 540
x"fdf60",-- -522
x"f8300",-- -2000
x"f7a10",-- -2143
x"fbc90",-- -1079
x"00cf0",-- 207
x"008c0",-- 140
x"faee0",-- -1298
x"f9ab0",-- -1621
x"fa4b0",-- -1461
x"fcbb0",-- -837
x"00570",-- 87
x"02910",-- 657
x"02ad0",-- 685
x"ff180",-- -232
x"ff4c0",-- -180
x"03bd0",-- 957
x"08000",-- 2048
x"0b8b0",-- 2955
x"0c230",-- 3107
x"0b010",-- 2817
x"0b360",-- 2870
x"0dd80",-- 3544
x"140c0",-- 5132
x"17e10",-- 6113
x"183e0",-- 6206
x"18910",-- 6289
x"175a0",-- 5978
x"18780",-- 6264
x"1b6f0",-- 7023
x"19a80",-- 6568
x"190f0",-- 6415
x"1e220",-- 7714
x"1ffb0",-- 8187
x"1ac80",-- 6856
x"11d70",-- 4567
x"110d0",-- 4365
x"17bf0",-- 6079
x"17a50",-- 6053
x"109b0",-- 4251
x"08d40",-- 2260
x"006e0",-- 110
x"fc520",-- -942
x"fffe0",-- -2
x"03590",-- 857
x"fa990",-- -1383
x"ec960",-- -4970
x"e8420",-- -6078
x"eb830",-- -5245
x"eda70",-- -4697
x"eb9f0",-- -5217
x"e9900",-- -5744
x"e5f10",-- -6671
x"e0190",-- -8167
x"e24b0",-- -7605
x"e9a20",-- -5726
x"e9f70",-- -5641
x"e66a0",-- -6550
x"e7770",-- -6281
x"e9fc0",-- -5636
x"e7ce0",-- -6194
x"e8120",-- -6126
x"eebc0",-- -4420
x"f34d0",-- -3251
x"f1c20",-- -3646
x"ef920",-- -4206
x"f0c50",-- -3899
x"f31a0",-- -3302
x"f57e0",-- -2690
x"fc160",-- -1002
x"febc0",-- -324
x"f8c80",-- -1848
x"f6070",-- -2553
x"fc430",-- -957
x"02190",-- 537
x"033b0",-- 827
x"03680",-- 872
x"02870",-- 647
x"00000",-- 0
x"ff170",-- -233
x"05c10",-- 1473
x"0c4b0",-- 3147
x"08e30",-- 2275
x"03d00",-- 976
x"02340",-- 564
x"03940",-- 916
x"06230",-- 1571
x"08370",-- 2103
x"085e0",-- 2142
x"02c10",-- 705
x"fb7b0",-- -1157
x"fa6c0",-- -1428
x"02f70",-- 759
x"059f0",-- 1439
x"00020",-- 2
x"fb240",-- -1244
x"f6190",-- -2535
x"f72f0",-- -2257
x"fdc70",-- -569
x"00bb0",-- 187
x"fd5b0",-- -677
x"f6960",-- -2410
x"f4990",-- -2919
x"f96d0",-- -1683
x"ff010",-- -255
x"ff990",-- -103
x"fcdf0",-- -801
x"fc480",-- -952
x"fb560",-- -1194
x"fddf0",-- -545
x"04850",-- 1157
x"075e0",-- 1886
x"06ed0",-- 1773
x"06760",-- 1654
x"07770",-- 1911
x"0af40",-- 2804
x"0ef40",-- 3828
x"13400",-- 4928
x"14110",-- 5137
x"137d0",-- 4989
x"146d0",-- 5229
x"17df0",-- 6111
x"1bee0",-- 7150
x"1d190",-- 7449
x"1e460",-- 7750
x"1bfd0",-- 7165
x"13bf0",-- 5055
x"17b50",-- 6069
x"23b40",-- 9140
x"238a0",-- 9098
x"1a6d0",-- 6765
x"0e0c0",-- 3596
x"0f8f0",-- 3983
x"16860",-- 5766
x"13e90",-- 5097
x"10410",-- 4161
x"08890",-- 2185
x"fc520",-- -942
x"f78b0",-- -2165
x"fdae0",-- -594
x"01060",-- 262
x"f5400",-- -2752
x"eafc0",-- -5380
x"ea170",-- -5609
x"e83c0",-- -6084
x"e72e0",-- -6354
x"e8280",-- -6104
x"ea600",-- -5536
x"e5ef0",-- -6673
x"de7b0",-- -8581
x"e1bb0",-- -7749
x"e68c0",-- -6516
x"e5810",-- -6783
x"e7470",-- -6329
x"eb950",-- -5227
x"e9d10",-- -5679
x"e3840",-- -7292
x"e7090",-- -6391
x"f1740",-- -3724
x"f4480",-- -3000
x"f2060",-- -3578
x"f0fc0",-- -3844
x"f1a90",-- -3671
x"f1de0",-- -3618
x"f7470",-- -2233
x"00a80",-- 168
x"ff1f0",-- -225
x"f8390",-- -1991
x"f9270",-- -1753
x"ff3b0",-- -197
x"02c60",-- 710
x"03fb0",-- 1019
x"05b50",-- 1461
x"04930",-- 1171
x"01770",-- 375
x"037b0",-- 891
x"085c0",-- 2140
x"07310",-- 1841
x"05ba0",-- 1466
x"08c00",-- 2240
x"08c00",-- 2240
x"04530",-- 1107
x"004e0",-- 78
x"038a0",-- 906
x"06390",-- 1593
x"03f80",-- 1016
x"01260",-- 294
x"fd920",-- -622
x"fb620",-- -1182
x"f8d50",-- -1835
x"fd800",-- -640
x"019a0",-- 410
x"f9740",-- -1676
x"f4d50",-- -2859
x"f6440",-- -2492
x"f7a10",-- -2143
x"fa610",-- -1439
x"fb7b0",-- -1157
x"fb390",-- -1223
x"f7d30",-- -2093
x"f6cd0",-- -2355
x"fb990",-- -1127
x"ff7b0",-- -133
x"00b70",-- 183
x"ff4e0",-- -178
x"00d20",-- 210
x"038b0",-- 907
x"040d0",-- 1037
x"08020",-- 2050
x"0c7c0",-- 3196
x"0cf20",-- 3314
x"0cd90",-- 3289
x"0f090",-- 3849
x"13790",-- 4985
x"14500",-- 5200
x"159b0",-- 5531
x"19640",-- 6500
x"1b3d0",-- 6973
x"1ba50",-- 7077
x"1bf10",-- 7153
x"1d670",-- 7527
x"1eac0",-- 7852
x"18340",-- 6196
x"15cb0",-- 5579
x"211c0",-- 8476
x"23690",-- 9065
x"1ab60",-- 6838
x"0eef0",-- 3823
x"0e890",-- 3721
x"15ff0",-- 5631
x"14180",-- 5144
x"0fe90",-- 4073
x"08250",-- 2085
x"fb830",-- -1149
x"f6de0",-- -2338
x"fc670",-- -921
x"01010",-- 257
x"f6fc0",-- -2308
x"e7c50",-- -6203
x"e5d60",-- -6698
x"e82e0",-- -6098
x"e7f20",-- -6158
x"e6c90",-- -6455
x"e75b0",-- -6309
x"e3890",-- -7287
x"dba00",-- -9312
x"dfdb0",-- -8229
x"e7ca0",-- -6198
x"e5a10",-- -6751
x"e3900",-- -7280
x"e7d40",-- -6188
x"e9f60",-- -5642
x"e5b30",-- -6733
x"e6d30",-- -6445
x"f0140",-- -4076
x"f3c90",-- -3127
x"f2300",-- -3536
x"f1e30",-- -3613
x"f3f80",-- -3080
x"f4a50",-- -2907
x"f7930",-- -2157
x"00250",-- 37
x"02550",-- 597
x"fb6a0",-- -1174
x"fa430",-- -1469
x"00eb0",-- 235
x"064e0",-- 1614
x"05d10",-- 1489
x"05600",-- 1376
x"07760",-- 1910
x"02c00",-- 704
x"02cf0",-- 719
x"0a0d0",-- 2573
x"0b770",-- 2935
x"08860",-- 2182
x"05240",-- 1316
x"05310",-- 1329
x"06440",-- 1604
x"03ec0",-- 1004
x"04490",-- 1097
x"05290",-- 1321
x"02c60",-- 710
x"fce90",-- -791
x"f99a0",-- -1638
x"fe850",-- -379
x"fcbe0",-- -834
x"fc890",-- -887
x"fca20",-- -862
x"f50e0",-- -2802
x"f3c70",-- -3129
x"f69b0",-- -2405
x"fb920",-- -1134
x"fbf90",-- -1031
x"f66c0",-- -2452
x"f4690",-- -2967
x"f5ac0",-- -2644
x"f9f60",-- -1546
x"fdb50",-- -587
x"fe4e0",-- -434
x"fd940",-- -620
x"fab60",-- -1354
x"fd770",-- -649
x"042d0",-- 1069
x"08000",-- 2048
x"08c30",-- 2243
x"08780",-- 2168
x"0a910",-- 2705
x"0ba10",-- 2977
x"0f1c0",-- 3868
x"151a0",-- 5402
x"16540",-- 5716
x"15080",-- 5384
x"15be0",-- 5566
x"17d20",-- 6098
x"1b100",-- 6928
x"1e9a0",-- 7834
x"1ede0",-- 7902
x"1f8d0",-- 8077
x"1db20",-- 7602
x"1af60",-- 6902
x"15d20",-- 5586
x"18720",-- 6258
x"24400",-- 9280
x"20f70",-- 8439
x"16f50",-- 5877
x"0b810",-- 2945
x"0a410",-- 2625
x"13b70",-- 5047
x"13180",-- 4888
x"0d2b0",-- 3371
x"029d0",-- 669
x"f4ca0",-- -2870
x"f1ed0",-- -3603
x"f8ee0",-- -1810
x"fe210",-- -479
x"f2d20",-- -3374
x"e3610",-- -7327
x"e1b60",-- -7754
x"e1c90",-- -7735
x"e37e0",-- -7298
x"e6f00",-- -6416
x"e65b0",-- -6565
x"df4d0",-- -8371
x"d92f0",-- -9937
x"dee10",-- -8479
x"e54d0",-- -6835
x"e5790",-- -6791
x"e68d0",-- -6515
x"e9430",-- -5821
x"e9950",-- -5739
x"e69c0",-- -6500
x"e8f80",-- -5896
x"f30e0",-- -3314
x"f78d0",-- -2163
x"f6850",-- -2427
x"f6aa0",-- -2390
x"f6be0",-- -2370
x"f6780",-- -2440
x"fbd60",-- -1066
x"063e0",-- 1598
x"07120",-- 1810
x"ffb80",-- -72
x"fe7a0",-- -390
x"026b0",-- 619
x"06af0",-- 1711
x"0abe0",-- 2750
x"0bd00",-- 3024
x"09220",-- 2338
x"03da0",-- 986
x"03dd0",-- 989
x"06b40",-- 1716
x"0a230",-- 2595
x"0cc70",-- 3271
x"07270",-- 1831
x"04580",-- 1112
x"ffe20",-- -30
x"fc8a0",-- -886
x"04a20",-- 1186
x"07310",-- 1841
x"00670",-- 103
x"f77f0",-- -2177
x"f41c0",-- -3044
x"f6940",-- -2412
x"fb240",-- -1244
x"fe7d0",-- -387
x"f8670",-- -1945
x"f1290",-- -3799
x"eff10",-- -4111
x"f2df0",-- -3361
x"fa070",-- -1529
x"fb0c0",-- -1268
x"f6a70",-- -2393
x"f4e40",-- -2844
x"f5790",-- -2695
x"f9d30",-- -1581
x"fde20",-- -542
x"00eb0",-- 235
x"01470",-- 327
x"ffa30",-- -93
x"01f90",-- 505
x"05830",-- 1411
x"09490",-- 2377
x"0d150",-- 3349
x"0fab0",-- 4011
x"10780",-- 4216
x"0f3b0",-- 3899
x"11ba0",-- 4538
x"16230",-- 5667
x"187d0",-- 6269
x"1bd80",-- 7128
x"19a00",-- 6560
x"18e10",-- 6369
x"1c6e0",-- 7278
x"1dcb0",-- 7627
x"205e0",-- 8286
x"22050",-- 8709
x"1ede0",-- 7902
x"1c3b0",-- 7227
x"161d0",-- 5661
x"13d70",-- 5079
x"1f1e0",-- 7966
x"21240",-- 8484
x"1a2f0",-- 6703
x"0c630",-- 3171
x"059a0",-- 1434
x"0cb30",-- 3251
x"0dc10",-- 3521
x"0c020",-- 3074
x"04e50",-- 1253
x"f5430",-- -2749
x"eca80",-- -4952
x"ef590",-- -4263
x"f6b90",-- -2375
x"f37e0",-- -3202
x"e5ca0",-- -6710
x"df020",-- -8446
x"dc190",-- -9191
x"dcd30",-- -9005
x"e1050",-- -7931
x"e4850",-- -7035
x"e1f60",-- -7690
x"da010",-- -9727
x"daf50",-- -9483
x"e1950",-- -7787
x"e40a0",-- -7158
x"e6170",-- -6633
x"eb160",-- -5354
x"ed970",-- -4713
x"ea3d0",-- -5571
x"e97a0",-- -5766
x"f1340",-- -3788
x"f8160",-- -2026
x"fb1a0",-- -1254
x"fd540",-- -684
x"fd270",-- -729
x"f9ec0",-- -1556
x"faeb0",-- -1301
x"04ca0",-- 1226
x"0bb80",-- 3000
x"093f0",-- 2367
x"04f20",-- 1266
x"03860",-- 902
x"03f30",-- 1011
x"080d0",-- 2061
x"0d600",-- 3424
x"0eef0",-- 3823
x"08890",-- 2185
x"00ed0",-- 237
x"033f0",-- 831
x"08e10",-- 2273
x"09dd0",-- 2525
x"074a0",-- 1866
x"03380",-- 824
x"fecb0",-- -309
x"fb2a0",-- -1238
x"fe7a0",-- -390
x"00f40",-- 244
x"fc230",-- -989
x"f9470",-- -1721
x"f5680",-- -2712
x"f6df0",-- -2337
x"f6620",-- -2462
x"f3240",-- -3292
x"f8440",-- -1980
x"f5a60",-- -2650
x"f3ec0",-- -3092
x"f5150",-- -2795
x"f3ef0",-- -3089
x"f5e20",-- -2590
x"f7560",-- -2218
x"fb6a0",-- -1174
x"fcf70",-- -777
x"fa1e0",-- -1506
x"fa580",-- -1448
x"fdd10",-- -559
x"03fd0",-- 1021
x"06860",-- 1670
x"06820",-- 1666
x"07d00",-- 2000
x"07a30",-- 1955
x"0b4c0",-- 2892
x"111d0",-- 4381
x"138a0",-- 5002
x"126d0",-- 4717
x"11800",-- 4480
x"14840",-- 5252
x"17800",-- 6016
x"18270",-- 6183
x"192b0",-- 6443
x"19170",-- 6423
x"199b0",-- 6555
x"1b380",-- 6968
x"1bec0",-- 7148
x"1d350",-- 7477
x"1c2f0",-- 7215
x"1c360",-- 7222
x"1b740",-- 7028
x"1a550",-- 6741
x"12a00",-- 4768
x"0f860",-- 3974
x"196f0",-- 6511
x"1ade0",-- 6878
x"14a40",-- 5284
x"09060",-- 2310
x"03100",-- 784
x"05d50",-- 1493
x"060f0",-- 1551
x"07040",-- 1796
x"008f0",-- 143
x"f1880",-- -3704
x"e8f30",-- -5901
x"ead90",-- -5415
x"f1b30",-- -3661
x"ef130",-- -4333
x"e3de0",-- -7202
x"de820",-- -8574
x"dbb30",-- -9293
x"db3b0",-- -9413
x"e07d0",-- -8067
x"e50a0",-- -6902
x"e22e0",-- -7634
x"dca00",-- -9056
x"e0060",-- -8186
x"e55e0",-- -6818
x"e6710",-- -6543
x"e9060",-- -5882
x"eed20",-- -4398
x"f17c0",-- -3716
x"f0b70",-- -3913
x"f17f0",-- -3713
x"f5d30",-- -2605
x"f9480",-- -1720
x"fca50",-- -859
x"021c0",-- 540
x"03c20",-- 962
x"00440",-- 68
x"fdfd0",-- -515
x"03f40",-- 1012
x"09680",-- 2408
x"0a340",-- 2612
x"094a0",-- 2378
x"06080",-- 1544
x"01fb0",-- 507
x"033f0",-- 831
x"09880",-- 2440
x"0bbd0",-- 3005
x"081c0",-- 2076
x"01680",-- 360
x"00f20",-- 242
x"01ee0",-- 494
x"02870",-- 647
x"02fe0",-- 766
x"00300",-- 48
x"fcb70",-- -841
x"f8e80",-- -1816
x"fa710",-- -1423
x"f8ee0",-- -1810
x"f7b80",-- -2120
x"f6d70",-- -2345
x"f8140",-- -2028
x"f8260",-- -2010
x"f3d40",-- -3116
x"f3650",-- -3227
x"f5100",-- -2800
x"f7830",-- -2173
x"f9fb0",-- -1541
x"fab90",-- -1351
x"f9240",-- -1756
x"f7390",-- -2247
x"f9590",-- -1703
x"fffb0",-- -5
x"02e00",-- 736
x"03880",-- 904
x"022d0",-- 557
x"03a80",-- 936
x"06460",-- 1606
x"09a10",-- 2465
x"0e040",-- 3588
x"0efc0",-- 3836
x"0e340",-- 3636
x"0e700",-- 3696
x"11790",-- 4473
x"127a0",-- 4730
x"13770",-- 4983
x"14750",-- 5237
x"14f40",-- 5364
x"156c0",-- 5484
x"133f0",-- 4927
x"11ee0",-- 4590
x"15450",-- 5445
x"16220",-- 5666
x"15af0",-- 5551
x"159e0",-- 5534
x"144d0",-- 5197
x"12f90",-- 4857
x"14480",-- 5192
x"15260",-- 5414
x"139b0",-- 5019
x"0e950",-- 3733
x"09290",-- 2345
x"0da60",-- 3494
x"11360",-- 4406
x"10e30",-- 4323
x"0aa20",-- 2722
x"038f0",-- 911
x"01bc0",-- 444
x"00b20",-- 178
x"01510",-- 337
x"00cd0",-- 205
x"f9a60",-- -1626
x"f0b40",-- -3916
x"edd90",-- -4647
x"ee8f0",-- -4465
x"ef740",-- -4236
x"ea580",-- -5544
x"e79d0",-- -6243
x"e61a0",-- -6630
x"e3190",-- -7399
x"e3b80",-- -7240
x"e6bf0",-- -6465
x"e7ab0",-- -6229
x"e6370",-- -6601
x"e88a0",-- -6006
x"ebe50",-- -5147
x"ed380",-- -4808
x"ebfc0",-- -5124
x"ef220",-- -4318
x"f2df0",-- -3361
x"f57e0",-- -2690
x"f74a0",-- -2230
x"f9700",-- -1680
x"fa080",-- -1528
x"f9a60",-- -1626
x"fca70",-- -857
x"01170",-- 279
x"027d0",-- 637
x"00af0",-- 175
x"00670",-- 103
x"00e30",-- 227
x"015b0",-- 347
x"01540",-- 340
x"02b60",-- 694
x"01600",-- 352
x"00a00",-- 160
x"00b90",-- 185
x"00570",-- 87
x"005d0",-- 93
x"ff090",-- -247
x"fe930",-- -365
x"febe0",-- -322
x"fedc0",-- -292
x"fc960",-- -874
x"fc260",-- -986
x"fc620",-- -926
x"faeb0",-- -1301
x"fb920",-- -1134
x"fc1e0",-- -994
x"fbc40",-- -1084
x"fb2c0",-- -1236
x"faa50",-- -1371
x"fbda0",-- -1062
x"fd9e0",-- -610
x"fce60",-- -794
x"ff2e0",-- -210
x"ffa60",-- -90
x"002f0",-- 47
x"01950",-- 405
x"02a00",-- 672
x"02520",-- 594
x"04500",-- 1104
x"069a0",-- 1690
x"06a00",-- 1696
x"08b30",-- 2227
x"070d0",-- 1805
x"06be0",-- 1726
x"0af70",-- 2807
x"07220",-- 1826
x"092b0",-- 2347
x"0e090",-- 3593
x"06760",-- 1654
x"09da0",-- 2522
x"0a750",-- 2677
x"05fb0",-- 1531
x"07830",-- 1923
x"07f30",-- 2035
x"08b30",-- 2227
x"066e0",-- 1646
x"03ab0",-- 939
x"05060",-- 1286
x"05440",-- 1348
x"051a0",-- 1306
x"027f0",-- 639
x"04d20",-- 1234
x"057b0",-- 1403
x"02ac0",-- 684
x"046e0",-- 1134
x"04640",-- 1124
x"03240",-- 804
x"05e90",-- 1513
x"06e80",-- 1768
x"04bb0",-- 1211
x"06170",-- 1559
x"06140",-- 1556
x"05590",-- 1369
x"068b0",-- 1675
x"07350",-- 1845
x"08520",-- 2130
x"09030",-- 2307
x"072b0",-- 1835
x"06200",-- 1568
x"05cb0",-- 1483
x"047d0",-- 1149
x"04200",-- 1056
x"03b50",-- 949
x"019c0",-- 412
x"00690",-- 105
x"ff1f0",-- -225
x"fd8f0",-- -625
x"fc620",-- -926
x"fb520",-- -1198
x"f9fb0",-- -1541
x"f95b0",-- -1701
x"f8fa0",-- -1798
x"f8750",-- -1931
x"f8460",-- -1978
x"f7d00",-- -2096
x"f7200",-- -2272
x"f7400",-- -2240
x"f84b0",-- -1973
x"f8140",-- -2028
x"f8d90",-- -1831
x"f8c10",-- -1855
x"f8480",-- -1976
x"f8c60",-- -1850
x"f8570",-- -1961
x"f8520",-- -1966
x"f8840",-- -1916
x"f8410",-- -1983
x"f7ab0",-- -2133
x"f7fb0",-- -2053
x"f7430",-- -2237
x"f6480",-- -2488
x"f75c0",-- -2212
x"f63c0",-- -2500
x"f4960",-- -2922
x"f79c0",-- -2148
x"f78b0",-- -2165
x"f4f00",-- -2832
x"f73e0",-- -2242
x"f7970",-- -2153
x"f68c0",-- -2420
x"f7ef0",-- -2065
x"f89d0",-- -1891
x"f8fd0",-- -1795
x"fa350",-- -1483
x"fb450",-- -1211
x"fb9e0",-- -1122
x"fc5d0",-- -931
x"fcd70",-- -809
x"fdcc0",-- -564
x"fed20",-- -302
x"ffbd0",-- -67
x"00460",-- 70
x"002b0",-- 43
x"01040",-- 260
x"019e0",-- 414
x"02550",-- 597
x"02f40",-- 756
x"03440",-- 836
x"037b0",-- 891
x"03b30",-- 947
x"05170",-- 1303
x"05ae0",-- 1454
x"05bc0",-- 1468
x"06a50",-- 1701
x"06b60",-- 1718
x"06c20",-- 1730
x"07740",-- 1908
x"076d0",-- 1901
x"07450",-- 1861
x"07830",-- 1923
x"075e0",-- 1886
x"076f0",-- 1903
x"07580",-- 1880
x"06fc0",-- 1788
x"06780",-- 1656
x"05f60",-- 1526
x"05bc0",-- 1468
x"05670",-- 1383
x"04e10",-- 1249
x"04340",-- 1076
x"03ab0",-- 939
x"032c0",-- 812
x"02890",-- 649
x"026e0",-- 622
x"01db0",-- 475
x"01940",-- 404
x"014e0",-- 334
x"00dc0",-- 220
x"00b20",-- 178
x"00490",-- 73
x"001e0",-- 30
x"00ac0",-- 172
x"00340",-- 52
x"00080",-- 8
x"00800",-- 128
x"00320",-- 50
x"00840",-- 132
x"00cb0",-- 203
x"01400",-- 320
x"01ec0",-- 492
x"027a0",-- 634
x"02670",-- 615
x"03560",-- 854
x"040f0",-- 1039
x"04a50",-- 1189
x"06000",-- 1536
x"06610",-- 1633
x"06d90",-- 1753
x"06fc0",-- 1788
x"06ca0",-- 1738
x"06a50",-- 1701
x"06ae0",-- 1710
x"06930",-- 1683
x"05860",-- 1414
x"053a0",-- 1338
x"03f40",-- 1012
x"02b40",-- 692
x"02120",-- 530
x"00840",-- 132
x"ff5e0",-- -162
x"fefc0",-- -260
x"fd1b0",-- -741
x"fca50",-- -859
x"fc3a0",-- -966
x"fac30",-- -1341
x"fb060",-- -1274
x"fa280",-- -1496
x"f9df0",-- -1569
x"f9940",-- -1644
x"f9450",-- -1723
x"f8ed0",-- -1811
x"f8c80",-- -1848
x"f8cb0",-- -1845
x"f8840",-- -1916
x"f8af0",-- -1873
x"f8750",-- -1931
x"f8700",-- -1936
x"f8520",-- -1966
x"f8480",-- -1976
x"f8200",-- -2016
x"f8670",-- -1945
x"f8530",-- -1965
x"f8530",-- -1965
x"f8ee0",-- -1810
x"f8a30",-- -1885
x"f8ca0",-- -1846
x"f9200",-- -1760
x"f94a0",-- -1718
x"f9ea0",-- -1558
x"fa620",-- -1438
x"fae30",-- -1309
x"fb390",-- -1223
x"fb470",-- -1209
x"fbec0",-- -1044
x"fc9e0",-- -866
x"fd900",-- -624
x"fdef0",-- -529
x"fe570",-- -425
x"fecf0",-- -305
x"ff6c0",-- -148
x"000a0",-- 10
x"00b10",-- 177
x"014f0",-- 335
x"01620",-- 354
x"02230",-- 547
x"02aa0",-- 682
x"034f0",-- 847
x"03b70",-- 951
x"03f80",-- 1016
x"04780",-- 1144
x"05040",-- 1284
x"05600",-- 1376
x"05a90",-- 1449
x"05ef0",-- 1519
x"05e20",-- 1506
x"06020",-- 1538
x"06530",-- 1619
x"06440",-- 1604
x"05ee0",-- 1518
x"05ba0",-- 1466
x"057b0",-- 1403
x"055e0",-- 1374
x"052b0",-- 1323
x"04cd0",-- 1229
x"04990",-- 1177
x"03fb0",-- 1019
x"038b0",-- 907
x"03970",-- 919
x"03380",-- 824
x"02980",-- 664
x"02490",-- 585
x"02160",-- 534
x"01ad0",-- 429
x"01800",-- 384
x"01580",-- 344
x"00f40",-- 244
x"00c80",-- 200
x"00730",-- 115
x"003c0",-- 60
x"002f0",-- 47
x"fffb0",-- -5
x"ffda0",-- -38
x"ff9a0",-- -102
x"ff970",-- -105
x"ff5b0",-- -165
x"ff2b0",-- -213
x"ff2b0",-- -213
x"ff2e0",-- -210
x"fef30",-- -269
x"fef20",-- -270
x"feda0",-- -294
x"fec50",-- -315
x"feb90",-- -327
x"febb0",-- -325
x"fecb0",-- -309
x"febc0",-- -324
x"fed00",-- -304
x"fee10",-- -287
x"fefd0",-- -259
x"ff110",-- -239
x"ff2e0",-- -210
x"ff4e0",-- -178
x"ffa90",-- -87
x"ffce0",-- -50
x"fffe0",-- -2
x"00550",-- 85
x"00670",-- 103
x"00910",-- 145
x"00f90",-- 249
x"00f00",-- 240
x"011c0",-- 284
x"01290",-- 297
x"011f0",-- 287
x"011d0",-- 285
x"00f50",-- 245
x"011d0",-- 285
x"00b20",-- 178
x"00b20",-- 178
x"00700",-- 112
x"00210",-- 33
x"003f0",-- 63
x"ffae0",-- -82
x"ffb50",-- -75
x"ff790",-- -135
x"ff3f0",-- -193
x"ff2b0",-- -213
x"fee40",-- -284
x"fed70",-- -297
x"fe960",-- -362
x"fe9b0",-- -357
x"fe7b0",-- -389
x"fe760",-- -394
x"fe570",-- -425
x"fe2d0",-- -467
x"fe020",-- -510
x"fde40",-- -540
x"fde00",-- -544
x"fdc10",-- -575
x"fdba0",-- -582
x"fd720",-- -654
x"fd3d0",-- -707
x"fd470",-- -697
x"fd250",-- -731
x"fd1a0",-- -742
x"fd180",-- -744
x"fd250",-- -731
x"fd290",-- -727
x"fd2e0",-- -722
x"fd590",-- -679
x"fd6c0",-- -660
x"fdb50",-- -587
x"fdf80",-- -520
x"fe300",-- -464
x"fe6c0",-- -404
x"fe990",-- -359
x"ff070",-- -249
x"ff680",-- -152
x"ffc60",-- -58
x"00160",-- 22
x"00480",-- 72
x"00850",-- 133
x"00f50",-- 245
x"01530",-- 339
x"018f0",-- 399
x"01d00",-- 464
x"01ec0",-- 492
x"02200",-- 544
x"02620",-- 610
x"02700",-- 624
x"02940",-- 660
x"02b60",-- 694
x"02ac0",-- 684
x"02d20",-- 722
x"02e50",-- 741
x"02cf0",-- 719
x"02d60",-- 726
x"02d40",-- 724
x"02b10",-- 689
x"02a30",-- 675
x"02b40",-- 692
x"02a80",-- 680
x"02990",-- 665
x"02800",-- 640
x"02550",-- 597
x"024b0",-- 587
x"02350",-- 565
x"02030",-- 515
x"01f90",-- 505
x"01d30",-- 467
x"01920",-- 402
x"01470",-- 327
x"01170",-- 279
x"00e40",-- 228
x"009d0",-- 157
x"00750",-- 117
x"00280",-- 40
x"ffd10",-- -47
x"ff740",-- -140
x"ff380",-- -200
x"ff070",-- -249
x"fec50",-- -315
x"fe9e0",-- -354
x"fe5a0",-- -422
x"fe1b0",-- -485
x"fdf60",-- -522
x"fdce0",-- -562
x"fdcb0",-- -565
x"fdae0",-- -594
x"fd880",-- -632
x"fd7c0",-- -644
x"fd790",-- -647
x"fd7b0",-- -645
x"fd850",-- -635
x"fda10",-- -607
x"fdab0",-- -597
x"fd8f0",-- -625
x"fdc90",-- -567
x"fe030",-- -509
x"fe140",-- -492
x"fe440",-- -444
x"fe570",-- -425
x"fe870",-- -377
x"fe9b0",-- -357
x"fec10",-- -319
x"ff070",-- -249
x"ff270",-- -217
x"ff420",-- -190
x"ff630",-- -157
x"ff830",-- -125
x"ffb50",-- -75
x"ffe70",-- -25
x"00050",-- 5
x"00280",-- 40
x"00350",-- 53
x"005a0",-- 90
x"00870",-- 135
x"00990",-- 153
x"00bc0",-- 188
x"00c00",-- 192
x"00d90",-- 217
x"00f50",-- 245
x"00f20",-- 242
x"01100",-- 272
x"010b0",-- 267
x"011c0",-- 284
x"011f0",-- 287
x"01180",-- 280
x"011f0",-- 287
x"01090",-- 265
x"00f50",-- 245
x"01080",-- 264
x"00ef0",-- 239
x"00d50",-- 213
x"00cb0",-- 203
x"00a80",-- 168
x"008f0",-- 143
x"008c0",-- 140
x"008a0",-- 138
x"00550",-- 85
x"005a0",-- 90
x"004e0",-- 78
x"00390",-- 57
x"004d0",-- 77
x"002b0",-- 43
x"00280",-- 40
x"00200",-- 32
x"fff30",-- -13
x"00140",-- 20
x"fffd0",-- -3
x"ffe50",-- -27
x"ffdb0",-- -37
x"ffc60",-- -58
x"ffd10",-- -47
x"ffb70",-- -73
x"ffc20",-- -62
x"ffa40",-- -92
x"ffad0",-- -83
x"ffa60",-- -90
x"ff950",-- -107
x"ffa80",-- -88
x"ff8a0",-- -118
x"ff940",-- -108
x"ffad0",-- -83
x"ffcb0",-- -53
x"ffc20",-- -62
x"ffd10",-- -47
x"ffdf0",-- -33
x"ffdd0",-- -35
x"fffe0",-- -2
x"fff40",-- -12
x"00000",-- 0
x"00110",-- 17
x"fff90",-- -7
x"00190",-- 25
x"00210",-- 33
x"000f0",-- 15
x"002f0",-- 47
x"00230",-- 35
x"001b0",-- 27
x"00190",-- 25
x"00120",-- 18
x"00030",-- 3
x"00000",-- 0
x"fff80",-- -8
x"ffee0",-- -18
x"ffea0",-- -22
x"ffe00",-- -32
x"ffcb0",-- -53
x"ffc60",-- -58
x"ffae0",-- -82
x"ffa60",-- -90
x"ff940",-- -108
x"ff6d0",-- -147
x"ff800",-- -128
x"ff8d0",-- -115
x"ff6d0",-- -147
x"ff540",-- -172
x"ff510",-- -175
x"ff380",-- -200
x"ff3b0",-- -197
x"ff4c0",-- -180
x"ff380",-- -200
x"ff1f0",-- -225
x"ff1d0",-- -227
x"ff1a0",-- -230
x"ff220",-- -222
x"ff240",-- -220
x"ff2e0",-- -210
x"ff2e0",-- -210
x"ff2b0",-- -213
x"ff2c0",-- -212
x"ff220",-- -222
x"ff2b0",-- -213
x"ff180",-- -232
x"ff1d0",-- -227
x"ff1f0",-- -225
x"ff210",-- -223
x"ff240",-- -220
x"ff240",-- -220
x"ff360",-- -202
x"ff5d0",-- -163
x"ff600",-- -160
x"ff760",-- -138
x"ff790",-- -135
x"ff790",-- -135
x"ffa30",-- -93
x"ffb20",-- -78
x"ffd00",-- -48
x"ffc70",-- -57
x"ffdb0",-- -37
x"fff80",-- -8
x"000f0",-- 15
x"00160",-- 22
x"002b0",-- 43
x"00390",-- 57
x"00230",-- 35
x"00370",-- 55
x"00440",-- 68
x"00640",-- 100
x"00660",-- 102
x"00710",-- 113
x"007b0",-- 123
x"007d0",-- 125
x"008c0",-- 140
x"007f0",-- 127
x"008c0",-- 140
x"00960",-- 150
x"00940",-- 148
x"00990",-- 153
x"009d0",-- 157
x"00940",-- 148
x"008f0",-- 143
x"00930",-- 147
x"008c0",-- 140
x"00800",-- 128
x"00850",-- 133
x"00760",-- 118
x"005d0",-- 93
x"00670",-- 103
x"00670",-- 103
x"005a0",-- 90
x"00500",-- 80
x"00500",-- 80
x"00430",-- 67
x"00430",-- 67
x"00320",-- 50
x"002f0",-- 47
x"002a0",-- 42
x"00210",-- 33
x"00030",-- 3
x"00050",-- 5
x"00020",-- 2
x"fff30",-- -13
x"ffec0",-- -20
x"ffe20",-- -30
x"ffdd0",-- -35
x"ffb20",-- -78
x"ffd10",-- -47
x"ffc10",-- -63
x"ffb30",-- -77
x"ffb20",-- -78
x"ffa40",-- -92
x"ffda0",-- -38
x"ffb20",-- -78
x"ffc20",-- -62
x"ffbf0",-- -65
x"ffa30",-- -93
x"ffce0",-- -50
x"ffa90",-- -87
x"ffc90",-- -55
x"ffbc0",-- -68
x"ffa60",-- -90
x"ffd10",-- -47
x"ffc90",-- -55
x"ffe70",-- -25
x"ffd10",-- -47
x"ffdb0",-- -37
x"ffe00",-- -32
x"ffdf0",-- -33
x"fffb0",-- -5
x"fff90",-- -7
x"fffe0",-- -2
x"ffe70",-- -25
x"00000",-- 0
x"00020",-- 2
x"00050",-- 5
x"00020",-- 2
x"00020",-- 2
x"00000",-- 0
x"fffb0",-- -5
x"00030",-- 3
x"00020",-- 2
x"00000",-- 0
x"fffe0",-- -2
x"fff90",-- -7
x"00020",-- 2
x"fff40",-- -12
x"fff10",-- -15
x"fff90",-- -7
x"fff10",-- -15
x"fff40",-- -12
x"ffea0",-- -22
x"ffe70",-- -25
x"ffdd0",-- -35
x"ffdf0",-- -33
x"ffe50",-- -27
x"ffdd0",-- -35
x"ffd30",-- -45
x"ffce0",-- -50
x"ffd00",-- -48
x"ffd10",-- -47
x"ffc90",-- -55
x"ffdd0",-- -35
x"ffce0",-- -50
x"ffc90",-- -55
x"ffd30",-- -45
x"ffd80",-- -40
x"ffe20",-- -30
x"ffd50",-- -43
x"ffe20",-- -30
x"ffe40",-- -28
x"ffdb0",-- -37
x"ffe20",-- -30
x"ffe90",-- -23
x"ffea0",-- -22
x"ffe40",-- -28
x"ffe20",-- -30
x"ffee0",-- -18
x"ffe50",-- -27
x"ffd60",-- -42
x"ffe50",-- -27
x"ffea0",-- -22
x"ffef0",-- -17
x"ffe00",-- -32
x"fff80",-- -8
x"00020",-- 2
x"00000",-- 0
x"000d0",-- 13
x"000f0",-- 15
x"00190",-- 25
x"00120",-- 18
x"00160",-- 22
x"001b0",-- 27
x"00210",-- 33
x"001e0",-- 30
x"00140",-- 20
x"001e0",-- 30
x"00230",-- 35
x"00210",-- 33
x"002b0",-- 43
x"002b0",-- 43
x"001c0",-- 28
x"00260",-- 38
x"00280",-- 40
x"00230",-- 35
x"001e0",-- 30
x"001b0",-- 27
x"001b0",-- 27
x"000c0",-- 12
x"00140",-- 20
x"000c0",-- 12
x"000f0",-- 15
x"000d0",-- 13
x"00050",-- 5
x"00000",-- 0
x"fffe0",-- -2
x"fffe0",-- -2
x"fff80",-- -8
x"fffe0",-- -2
x"fffb0",-- -5
x"fff10",-- -15
x"ffe20",-- -30
x"ffdd0",-- -35
x"ffe20",-- -30
x"ffe20",-- -30
x"ffe50",-- -27
x"ffd50",-- -43
x"ffc70",-- -57
x"ffce0",-- -50
x"ffdb0",-- -37
x"ffe50",-- -27
x"ffd60",-- -42
x"ffdb0",-- -37
x"ffbd0",-- -67
x"ffce0",-- -50
x"ff9e0",-- -98
x"ffc40",-- -60
x"ff630",-- -157
x"ff740",-- -140
x"fe8c0",-- -372
x"fea20",-- -350
x"f9a80",-- -1624
x"f40f0",-- -3057
x"00480",-- 72
x"07e40",-- 2020
x"01810",-- 385
x"00760",-- 118
x"00870",-- 135
x"ff360",-- -202
x"02370",-- 567
x"01f10",-- 497
x"00480",-- 72
x"ff630",-- -157
x"fffe0",-- -2
x"019a0",-- 410
x"00cf0",-- 207
x"021c0",-- 540
x"03ab0",-- 939
x"02730",-- 627
x"02110",-- 529
x"01e70",-- 487
x"fff40",-- -12
x"ffbc0",-- -68
x"002a0",-- 42
x"005a0",-- 90
x"ff7c0",-- -132
x"ff740",-- -140
x"fed90",-- -295
x"ff110",-- -239
x"00980",-- 152
x"ff1f0",-- -225
x"ff040",-- -252
x"ffbf0",-- -65
x"ffe70",-- -25
x"ff8a0",-- -118
x"019e0",-- 414
x"01e20",-- 482
x"ff240",-- -220
x"00a70",-- 167
x"00440",-- 68
x"ff420",-- -190
x"03670",-- 871
x"00b90",-- 185
x"ff990",-- -103
x"02750",-- 629
x"ffc60",-- -58
x"01b20",-- 434
x"fb2c0",-- -1236
x"f1830",-- -3709
x"ffea0",-- -22
x"06390",-- 1593
x"f5680",-- -2712
x"f6480",-- -2488
x"03e90",-- 1001
x"02c50",-- 709
x"ff1d0",-- -227
x"ff060",-- -250
x"fdf90",-- -519
x"ffa60",-- -90
x"044b0",-- 1099
x"004b0",-- 75
x"fbf10",-- -1039
x"00de0",-- 222
x"04a00",-- 1184
x"024b0",-- 587
x"02c10",-- 705
x"02d70",-- 727
x"03010",-- 769
x"07220",-- 1826
x"01ce0",-- 462
x"00300",-- 48
x"06a70",-- 1703
x"ff810",-- -127
x"fd850",-- -635
x"03a40",-- 932
x"ffba0",-- -70
x"fc490",-- -951
x"02aa0",-- 682
x"fe0a0",-- -502
x"fe300",-- -464
x"ffee0",-- -18
x"feb20",-- -334
x"01770",-- 375
x"fe110",-- -495
x"fdfd0",-- -515
x"01970",-- 407
x"ff9c0",-- -100
x"fdfd0",-- -515
x"fd760",-- -650
x"fda80",-- -600
x"f9330",-- -1741
x"f8a00",-- -1888
x"00280",-- 40
x"fe870",-- -377
x"ff650",-- -155
x"fc610",-- -927
x"fd6f0",-- -657
x"ff3b0",-- -197
x"011a0",-- 282
x"05fe0",-- 1534
x"01ad0",-- 429
x"fe2d0",-- -467
x"03a80",-- 936
x"048c0",-- 1164
x"ff740",-- -140
x"00610",-- 97
x"07350",-- 1845
x"02aa0",-- 682
x"033a0",-- 826
x"051a0",-- 1306
x"02a20",-- 674
x"00eb0",-- 235
x"01060",-- 262
x"04670",-- 1127
x"fecf0",-- -305
x"ff350",-- -203
x"014a0",-- 330
x"fb390",-- -1223
x"fea00",-- -352
x"ffad0",-- -83
x"fceb0",-- -789
x"fdc70",-- -569
x"fafc0",-- -1284
x"febb0",-- -325
x"00ca0",-- 202
x"fe750",-- -395
x"ff420",-- -190
x"fa140",-- -1516
x"01290",-- 297
x"fe3a0",-- -454
x"fd420",-- -702
x"02550",-- 597
x"f8cb0",-- -1845
x"02670",-- 615
x"00c60",-- 198
x"fdb80",-- -584
x"05bc0",-- 1468
x"ff510",-- -175
x"02e30",-- 739
x"05cb0",-- 1483
x"fe020",-- -510
x"054c0",-- 1356
x"00960",-- 150
x"ff110",-- -239
x"02ad0",-- 685
x"ff0c0",-- -244
x"05760",-- 1398
x"ff310",-- -207
x"02bc0",-- 700
x"03cb0",-- 971
x"00120",-- 18
x"00250",-- 37
x"034f0",-- 847
x"fe140",-- -492
x"fe300",-- -464
x"05400",-- 1344
x"fa0c0",-- -1524
x"03300",-- 816
x"fca70",-- -857
x"01710",-- 369
x"ff4e0",-- -178
x"00cd0",-- 205
x"01a90",-- 425
x"ff270",-- -217
x"00a00",-- 160
x"ff2c0",-- -212
x"00f70",-- 247
x"fb740",-- -1164
x"060d0",-- 1549
x"fb670",-- -1177
x"fd590",-- -679
x"03e50",-- 997
x"f9c40",-- -1596
x"fcb60",-- -842
x"fb240",-- -1244
x"fc990",-- -871
x"04200",-- 1056
x"fd9c0",-- -612
x"fe1e0",-- -482
x"07ef0",-- 2031
x"fac80",-- -1336
x"016a0",-- 362
x"01ab0",-- 427
x"fb250",-- -1243
x"02260",-- 550
x"fd340",-- -716
x"04500",-- 1104
x"00d00",-- 208
x"f7970",-- -2153
x"08980",-- 2200
x"02c30",-- 707
x"f9b20",-- -1614
x"07170",-- 1815
x"03680",-- 872
x"fbc40",-- -1084
x"00df0",-- 223
x"02370",-- 567
x"f91d0",-- -1763
x"08770",-- 2167
x"fc5c0",-- -932
x"fc660",-- -922
x"06750",-- 1653
x"fdb20",-- -590
x"fcd00",-- -816
x"fdfd0",-- -515
x"04ae0",-- 1198
x"faca0",-- -1334
x"ff2e0",-- -210
x"05530",-- 1363
x"fd100",-- -752
x"01900",-- 400
x"01c20",-- 450
x"f9b50",-- -1611
x"04b10",-- 1201
x"fd9a0",-- -614
x"fba40",-- -1116
x"06f50",-- 1781
x"fce10",-- -799
x"fe930",-- -365
x"04390",-- 1081
x"f8f50",-- -1803
x"019e0",-- 414
x"06c50",-- 1733
x"f8190",-- -2023
x"058f0",-- 1423
x"03cc0",-- 972
x"f8b20",-- -1870
x"02e10",-- 737
x"00350",-- 53
x"fdfd0",-- -515
x"fe3e0",-- -450
x"023f0",-- 575
x"00dc0",-- 220
x"fd9c0",-- -612
x"006b0",-- 107
x"fec80",-- -312
x"fba80",-- -1112
x"fed70",-- -297
x"fa940",-- -1388
x"00c10",-- 193
x"00bc0",-- 188
x"faa00",-- -1376
x"fc1c0",-- -996
x"01b50",-- 437
x"fd160",-- -746
x"03420",-- 834
x"010d0",-- 269
x"fd600",-- -672
x"05120",-- 1298
x"ff350",-- -203
x"033b0",-- 827
x"02870",-- 647
x"ffa60",-- -90
x"02660",-- 614
x"05fd0",-- 1533
x"049d0",-- 1181
x"fcc00",-- -832
x"042d0",-- 1069
x"fe190",-- -487
x"02b20",-- 690
x"01880",-- 392
x"02340",-- 564
x"015e0",-- 350
x"f9240",-- -1756
x"028a0",-- 650
x"ffec0",-- -20
x"fc910",-- -879
x"fefd0",-- -259
x"009d0",-- 157
x"f8640",-- -1948
x"fff40",-- -12
x"053b0",-- 1339
x"fa250",-- -1499
x"fe410",-- -447
x"02430",-- 579
x"fdc70",-- -569
x"007d0",-- 125
x"06250",-- 1573
x"fb250",-- -1243
x"fcbb0",-- -837
x"06570",-- 1623
x"fda40",-- -604
x"ffa30",-- -93
x"04350",-- 1077
x"fe390",-- -455
x"fe2b0",-- -469
x"04a50",-- 1189
x"ffa30",-- -93
x"00dc0",-- 220
x"02840",-- 644
x"fceb0",-- -789
x"028a0",-- 650
x"ffc20",-- -62
x"01c60",-- 454
x"01260",-- 294
x"fd2e0",-- -722
x"01710",-- 369
x"011c0",-- 284
x"ffce0",-- -50
x"f9330",-- -1741
x"05d10",-- 1489
x"feaa0",-- -342
x"f7630",-- -2205
x"0a780",-- 2680
x"fcaa0",-- -854
x"f95e0",-- -1698
x"06e60",-- 1766
x"fa9d0",-- -1379
x"ff400",-- -192
x"04d10",-- 1233
x"ff3d0",-- -195
x"fd330",-- -717
x"00500",-- 80
x"01e90",-- 489
x"fde50",-- -539
x"00350",-- 53
x"ff3a0",-- -198
x"03090",-- 777
x"fd1d0",-- -739
x"ff510",-- -175
x"04eb0",-- 1259
x"fb420",-- -1214
x"ffb20",-- -78
x"04910",-- 1169
x"fe7f0",-- -385
x"fc050",-- -1019
x"06e30",-- 1763
x"00750",-- 117
x"f9a40",-- -1628
x"01940",-- 404
x"02f90",-- 761
x"fde90",-- -535
x"fed70",-- -297
x"03a40",-- 932
x"fdb70",-- -585
x"013d0",-- 317
x"01150",-- 277
x"fcf00",-- -784
x"02ed0",-- 749
x"00f20",-- 242
x"fc430",-- -957
x"02840",-- 644
x"00200",-- 32
x"fef30",-- -269
x"010d0",-- 269
x"ffe40",-- -28
x"fccd0",-- -819
x"052b0",-- 1323
x"ff2e0",-- -210
x"fa6e0",-- -1426
x"062d0",-- 1581
x"fa020",-- -1534
x"fe070",-- -505
x"06aa0",-- 1706
x"f9540",-- -1708
x"fbef0",-- -1041
x"07860",-- 1926
x"fb850",-- -1147
x"fd680",-- -664
x"00c10",-- 193
x"01ce0",-- 462
x"010b0",-- 267
x"fc5c0",-- -932
x"00030",-- 3
x"02fc0",-- 764
x"fe0c0",-- -500
x"fe0a0",-- -502
x"03b30",-- 947
x"fecf0",-- -305
x"00230",-- 35
x"047b0",-- 1147
x"fe1e0",-- -482
x"fdab0",-- -597
x"07670",-- 1895
x"f9560",-- -1706
x"ffbd0",-- -67
x"05490",-- 1353
x"fb710",-- -1167
x"00a00",-- 160
x"00280",-- 40
x"feb20",-- -334
x"fbe00",-- -1056
x"03c40",-- 964
x"012c0",-- 300
x"f7d80",-- -2088
x"0a2d0",-- 2605
x"fda40",-- -604
x"f8190",-- -2023
x"09450",-- 2373
x"faad0",-- -1363
x"feb40",-- -332
x"035e0",-- 862
x"fdb20",-- -590
x"03920",-- 914
x"f9990",-- -1639
x"018d0",-- 397
x"05ea0",-- 1514
x"f8960",-- -1898
x"02e00",-- 736
x"03990",-- 921
x"fdfd0",-- -515
x"02350",-- 565
x"ffa60",-- -90
x"fcb20",-- -846
x"03420",-- 834
x"00250",-- 37
x"fb310",-- -1231
x"05130",-- 1299
x"fccd0",-- -819
x"fbe40",-- -1052
x"03590",-- 857
x"00ed0",-- 237
x"ff9a0",-- -102
x"fee80",-- -280
x"00320",-- 50
x"01490",-- 329
x"00110",-- 17
x"fa190",-- -1511
x"03e40",-- 996
x"040a0",-- 1034
x"f6a20",-- -2398
x"042d0",-- 1069
x"080f0",-- 2063
x"f6370",-- -2505
x"00f50",-- 245
x"05ce0",-- 1486
x"fafd0",-- -1283
x"02e10",-- 737
x"00760",-- 118
x"f8730",-- -1933
x"02be0",-- 702
x"06490",-- 1609
x"f80d0",-- -2035
x"03130",-- 787
x"05940",-- 1428
x"f7090",-- -2295
x"05010",-- 1281
x"00c80",-- 200
x"fd200",-- -736
x"025a0",-- 602
x"fd880",-- -632
x"fcda0",-- -806
x"03bd0",-- 957
x"06e60",-- 1766
x"f91b0",-- -1765
x"fe030",-- -509
x"05dd0",-- 1501
x"fc340",-- -972
x"008c0",-- 140
x"060a0",-- 1546
x"f8e60",-- -1818
x"02dc0",-- 732
x"02800",-- 640
x"fe320",-- -462
x"04170",-- 1047
x"fa780",-- -1416
x"00120",-- 18
x"046c0",-- 1132
x"fd880",-- -632
x"043e0",-- 1086
x"fdd80",-- -552
x"fe700",-- -400
x"01940",-- 404
x"fdf30",-- -525
x"05530",-- 1363
x"febb0",-- -325
x"fe250",-- -475
x"fcb60",-- -842
x"024b0",-- 587
x"000d0",-- 13
x"fa170",-- -1513
x"002b0",-- 43
x"036f0",-- 879
x"fcc50",-- -827
x"f7400",-- -2240
x"06570",-- 1623
x"fcc80",-- -824
x"ffb80",-- -72
x"fd620",-- -670
x"ff220",-- -222
x"092e0",-- 2350
x"fa710",-- -1423
x"01e50",-- 485
x"fe960",-- -362
x"00250",-- 37
x"062b0",-- 1579
x"fd800",-- -640
x"03da0",-- 986
x"03c70",-- 967
x"fd1b0",-- -741
x"060f0",-- 1551
x"fc580",-- -936
x"02140",-- 532
x"07e00",-- 2016
x"fa730",-- -1421
x"ff950",-- -107
x"08140",-- 2068
x"ff210",-- -223
x"fa050",-- -1531
x"02340",-- 564
x"feda0",-- -294
x"007d0",-- 125
x"026b0",-- 619
x"fc580",-- -936
x"01f90",-- 505
x"03a40",-- 932
x"f9b80",-- -1608
x"03130",-- 787
x"03b80",-- 952
x"fe430",-- -445
x"00050",-- 5
x"027f0",-- 639
x"02ad0",-- 685
x"fd1a0",-- -742
x"003e0",-- 62
x"033d0",-- 829
x"034f0",-- 847
x"fb7e0",-- -1154
x"049e0",-- 1182
x"04080",-- 1032
x"fd020",-- -766
x"ff2b0",-- -213
x"018d0",-- 397
x"030d0",-- 781
x"fae60",-- -1306
x"04140",-- 1044
x"06340",-- 1588
x"fcb40",-- -844
x"f98a0",-- -1654
x"011c0",-- 284
x"05350",-- 1333
x"fd290",-- -727
x"fdd60",-- -554
x"01c20",-- 450
x"ff510",-- -175
x"ffa90",-- -87
x"fceb0",-- -789
x"024e0",-- 590
x"03bd0",-- 957
x"f7720",-- -2190
x"ff950",-- -107
x"086e0",-- 2158
x"fea00",-- -352
x"fc500",-- -944
x"02bb0",-- 699
x"00050",-- 5
x"00570",-- 87
x"02b90",-- 697
x"01cb0",-- 459
x"02a30",-- 675
x"fbd10",-- -1071
x"fd290",-- -727
x"09150",-- 2325
x"fe0a0",-- -502
x"fd100",-- -752
x"03b00",-- 944
x"fb0b0",-- -1269
x"02200",-- 544
x"01010",-- 257
x"fc0c0",-- -1012
x"02bc0",-- 700
x"fd4c0",-- -692
x"fe6e0",-- -402
x"05ad0",-- 1453
x"fdea0",-- -534
x"fd600",-- -672
x"fe5c0",-- -420
x"021c0",-- 540
x"02f40",-- 756
x"ff8d0",-- -115
x"fd1a0",-- -742
x"feb40",-- -332
x"ff290",-- -215
x"ff070",-- -249
x"05b20",-- 1458
x"fcc30",-- -829
x"ff220",-- -222
x"02980",-- 664
x"f7d80",-- -2088
x"06480",-- 1608
x"04230",-- 1059
x"f62a0",-- -2518
x"07330",-- 1843
x"01ef0",-- 495
x"f90b0",-- -1781
x"020d0",-- 525
x"02940",-- 660
x"f9970",-- -1641
x"06210",-- 1569
x"02fa0",-- 762
x"f41c0",-- -3044
x"03d10",-- 977
x"085f0",-- 2143
x"fbf30",-- -1037
x"fe0a0",-- -502
x"019e0",-- 414
x"fcbb0",-- -837
x"035d0",-- 861
x"ff150",-- -235
x"fe9b0",-- -357
x"04aa0",-- 1194
x"f85d0",-- -1955
x"fc520",-- -942
x"0e8c0",-- 3724
x"f9bc0",-- -1604
x"f3130",-- -3309
x"0a860",-- 2694
x"fdb80",-- -584
x"fb6c0",-- -1172
x"07260",-- 1830
x"fa0f0",-- -1521
x"fa640",-- -1436
x"065d0",-- 1629
x"fecd0",-- -307
x"05c70",-- 1479
x"00000",-- 0
x"f2d70",-- -3369
x"050b0",-- 1291
x"06460",-- 1606
x"fe210",-- -479
x"fde40",-- -540
x"03c10",-- 961
x"027f0",-- 639
x"f8960",-- -1898
x"00070",-- 7
x"08ed0",-- 2285
x"ff9f0",-- -97
x"f89e0",-- -1890
x"02ff0",-- 767
x"05e20",-- 1506
x"ff620",-- -158
x"f95b0",-- -1701
x"fd160",-- -746
x"065c0",-- 1628
x"fe500",-- -432
x"fb3d0",-- -1219
x"04520",-- 1106
x"feda0",-- -294
x"fa8a0",-- -1398
x"01010",-- 257
x"04a20",-- 1186
x"00230",-- 35
x"f73b0",-- -2245
x"02b70",-- 695
x"07380",-- 1848
x"f8940",-- -1900
x"fc660",-- -922
x"08230",-- 2083
x"000d0",-- 13
x"f8030",-- -2045
x"01a30",-- 419
x"07a30",-- 1955
x"fc660",-- -922
x"f84b0",-- -1973
x"05a30",-- 1443
x"04be0",-- 1214
x"fe3e0",-- -450
x"fc350",-- -971
x"fee10",-- -287
x"06870",-- 1671
x"fa6c0",-- -1428
x"fb990",-- -1127
x"07c70",-- 1991
x"00a20",-- 162
x"f59c0",-- -2660
x"00700",-- 112
x"08b60",-- 2230
x"fe750",-- -395
x"fc6e0",-- -914
x"fbfd0",-- -1027
x"019a0",-- 410
x"03bc0",-- 956
x"faf70",-- -1289
x"01900",-- 400
x"09170",-- 2327
x"f7400",-- -2240
x"f7130",-- -2285
x"0c8b0",-- 3211
x"05800",-- 1408
x"f5090",-- -2807
x"042a0",-- 1066
x"03510",-- 849
x"f94a0",-- -1718
x"010e0",-- 270
x"003e0",-- 62
x"ff830",-- -125
x"02a30",-- 675
x"ffee0",-- -18
x"ffe90",-- -23
x"02aa0",-- 682
x"fc730",-- -909
x"fc8e0",-- -882
x"016d0",-- 365
x"04250",-- 1061
x"fe3a0",-- -454
x"fbec0",-- -1044
x"03760",-- 886
x"022a0",-- 554
x"f93e0",-- -1730
x"01240",-- 292
x"094c0",-- 2380
x"fe760",-- -394
x"f8de0",-- -1826
x"033f0",-- 831
x"04b40",-- 1204
x"f83a0",-- -1990
x"02200",-- 544
x"04cf0",-- 1231
x"fb9f0",-- -1121
x"00410",-- 65
x"fd720",-- -654
x"02430",-- 579
x"05ab0",-- 1451
x"f8e30",-- -1821
x"ff880",-- -120
x"030b0",-- 779
x"fa0a0",-- -1526
x"ff440",-- -188
x"04550",-- 1109
x"fe460",-- -442
x"fe200",-- -480
x"ffd80",-- -40
x"fea00",-- -352
x"06440",-- 1604
x"fd1a0",-- -742
x"f7400",-- -2240
x"09bd0",-- 2493
x"03e00",-- 992
x"f6de0",-- -2338
x"03580",-- 856
x"04490",-- 1097
x"fb160",-- -1258
x"03cc0",-- 972
x"03c60",-- 966
x"fcb20",-- -846
x"fff80",-- -8
x"fcbe0",-- -834
x"ff070",-- -249
x"074a0",-- 1866
x"015e0",-- 350
x"feb20",-- -334
x"01e70",-- 487
x"fc6c0",-- -916
x"000c0",-- 12
x"01df0",-- 479
x"fc3c0",-- -964
x"ff240",-- -220
x"ff8a0",-- -118
x"00ad0",-- 173
x"01e90",-- 489
x"ffbf0",-- -65
x"fed40",-- -300
x"fced0",-- -787
x"ff760",-- -138
x"027b0",-- 635
x"02430",-- 579
x"fd470",-- -697
x"006e0",-- 110
x"010d0",-- 269
x"005f0",-- 95
x"04a90",-- 1193
x"ff790",-- -135
x"fd8f0",-- -625
x"fec50",-- -315
x"035e0",-- 862
x"011d0",-- 285
x"00760",-- 118
x"03720",-- 882
x"fab90",-- -1351
x"fd420",-- -702
x"05620",-- 1378
x"02e80",-- 744
x"fd8d0",-- -627
x"ff440",-- -188
x"ff0c0",-- -244
x"fd860",-- -634
x"ff090",-- -247
x"febc0",-- -324
x"00f90",-- 249
x"fe440",-- -444
x"02f20",-- 754
x"00840",-- 132
x"f9a30",-- -1629
x"00e10",-- 225
x"fe9b0",-- -357
x"fc6c0",-- -916
x"05100",-- 1296
x"040c0",-- 1036
x"fe000",-- -512
x"fd020",-- -766
x"ff8b0",-- -117
x"02500",-- 592
x"fdc20",-- -574
x"ff580",-- -168
x"030d0",-- 781
x"00c00",-- 192
x"fead0",-- -339
x"02990",-- 665
x"fd830",-- -637
x"fddf0",-- -545
x"03ba0",-- 954
x"fd110",-- -751
x"015b0",-- 347
x"024b0",-- 587
x"fe1b0",-- -485
x"00430",-- 67
x"fc9e0",-- -866
x"ffe20",-- -30
x"ffd50",-- -43
x"fc6e0",-- -914
x"00800",-- 128
x"02190",-- 537
x"ffb70",-- -73
x"fbea0",-- -1046
x"fe7f0",-- -385
x"ff760",-- -138
x"fe6b0",-- -405
x"ff5b0",-- -165
x"fe460",-- -442
x"00350",-- 53
x"00530",-- 83
x"fe3e0",-- -450
x"fdfb0",-- -517
x"01a90",-- 425
x"fe9b0",-- -357
x"fc780",-- -904
x"06c50",-- 1733
x"03a90",-- 937
x"fa170",-- -1513
x"fce40",-- -796
x"00d20",-- 210
x"01490",-- 329
x"fe6c0",-- -404
x"ff380",-- -200
x"043c0",-- 1084
x"ff540",-- -172
x"faaa0",-- -1366
x"03450",-- 837
x"02aa0",-- 682
x"fd2c0",-- -724
x"fd650",-- -667
x"019f0",-- 415
x"02890",-- 649
x"fe960",-- -362
x"01fd0",-- 509
x"fdee0",-- -530
x"ff970",-- -105
x"04620",-- 1122
x"fc7d0",-- -899
x"fe190",-- -487
x"04530",-- 1107
x"fdda0",-- -550
x"ff470",-- -185
x"05580",-- 1368
x"ff020",-- -254
x"fe030",-- -509
x"00480",-- 72
x"015e0",-- 350
x"ff600",-- -160
x"fef30",-- -269
x"03ab0",-- 939
x"ff260",-- -218
x"fb650",-- -1179
x"03150",-- 789
x"03120",-- 786
x"ff540",-- -172
x"021c0",-- 540
x"00250",-- 37
x"fdd10",-- -559
x"02cf0",-- 719
x"008f0",-- 143
x"fddd0",-- -547
x"02fe0",-- 766
x"04cd0",-- 1229
x"ff510",-- -175
x"fdf10",-- -527
x"06eb0",-- 1771
x"006c0",-- 108
x"fcc80",-- -824
x"05c20",-- 1474
x"04030",-- 1027
x"ffda0",-- -38
x"00840",-- 132
x"031d0",-- 797
x"00f00",-- 240
x"fec60",-- -314
x"047f0",-- 1151
x"056c0",-- 1388
x"fe7b0",-- -389
x"fe3a0",-- -454
x"03cc0",-- 972
x"02370",-- 567
x"fdd10",-- -559
x"00780",-- 120
x"038f0",-- 911
x"00280",-- 40
x"fe580",-- -424
x"01ad0",-- 429
x"017b0",-- 379
x"fec80",-- -312
x"ffcc0",-- -52
x"ffc90",-- -55
x"ffc40",-- -60
x"ffb00",-- -80
x"ff680",-- -152
x"01710",-- 369
x"00e40",-- 228
x"ffc90",-- -55
x"002a0",-- 42
x"ff220",-- -222
x"fe140",-- -492
x"ffea0",-- -22
x"00050",-- 5
x"000f0",-- 15
x"fda30",-- -605
x"fc580",-- -936
x"ff270",-- -217
x"fe050",-- -507
x"fccd0",-- -819
x"fd590",-- -679
x"ff3a0",-- -198
x"fd2a0",-- -726
x"f9160",-- -1770
x"fd360",-- -714
x"fd8b0",-- -629
x"fa710",-- -1423
x"fc8e0",-- -882
x"fdae0",-- -594
x"fb6c0",-- -1172
x"f8c50",-- -1851
x"fa3f0",-- -1473
x"fe070",-- -505
x"fb710",-- -1167
x"fa300",-- -1488
x"fd2e0",-- -722
x"fe030",-- -509
x"fabc0",-- -1348
x"fa2b0",-- -1493
x"fec80",-- -312
x"fe530",-- -429
x"fa000",-- -1536
x"f9da0",-- -1574
x"fff80",-- -8
x"00f00",-- 240
x"f8c00",-- -1856
x"fba90",-- -1111
x"03470",-- 839
x"fe480",-- -440
x"faa00",-- -1376
x"ff670",-- -153
x"039c0",-- 924
x"ffb80",-- -72
x"fb880",-- -1144
x"00490",-- 73
x"04c70",-- 1223
x"fe4d0",-- -435
x"ff270",-- -217
x"04940",-- 1172
x"017e0",-- 382
x"fe9e0",-- -354
x"01a30",-- 419
x"0a950",-- 2709
x"036c0",-- 876
x"fe3e0",-- -450
x"0a6b0",-- 2667
x"0b1c0",-- 2844
x"fdf80",-- -520
x"02ca0",-- 714
x"0fc40",-- 4036
x"066c0",-- 1644
x"00d40",-- 212
x"0b150",-- 2837
x"0c930",-- 3219
x"070d0",-- 1805
x"05c90",-- 1481
x"06bb0",-- 1723
x"08e60",-- 2278
x"09c20",-- 2498
x"091f0",-- 2335
x"0d3b0",-- 3387
x"0d9a0",-- 3482
x"05270",-- 1319
x"04070",-- 1031
x"0b0b0",-- 2827
x"0ab60",-- 2742
x"06670",-- 1639
x"07e00",-- 2016
x"0dc90",-- 3529
x"09f40",-- 2548
x"01f40",-- 500
x"09a80",-- 2472
x"0e410",-- 3649
x"04f00",-- 1264
x"027d0",-- 637
x"0a2d0",-- 2605
x"07770",-- 1911
x"007d0",-- 125
x"024e0",-- 590
x"04e80",-- 1256
x"01440",-- 324
x"fb650",-- -1179
x"fc320",-- -974
x"fe460",-- -442
x"fa210",-- -1503
x"f5740",-- -2700
x"f8670",-- -1945
x"f7750",-- -2187
x"f0fa0",-- -3846
x"f2200",-- -3552
x"f5340",-- -2764
x"f28e0",-- -3442
x"ef830",-- -4221
x"ef1f0",-- -4321
x"f0530",-- -4013
x"f0af0",-- -3921
x"ee940",-- -4460
x"efd30",-- -4141
x"f2870",-- -3449
x"f0260",-- -4058
x"ef3e0",-- -4290
x"f2d70",-- -3369
x"f50e0",-- -2802
x"f2f30",-- -3341
x"f2990",-- -3431
x"f5720",-- -2702
x"f5da0",-- -2598
x"f5390",-- -2759
x"f8260",-- -2010
x"f87b0",-- -1925
x"f7220",-- -2270
x"f7600",-- -2208
x"f8850",-- -1915
x"fa580",-- -1448
x"fa350",-- -1483
x"f8fd0",-- -1795
x"fa2f0",-- -1489
x"fa5d0",-- -1443
x"fb150",-- -1259
x"fc230",-- -989
x"fbad0",-- -1107
x"fb430",-- -1213
x"faf00",-- -1296
x"ff650",-- -155
x"fdbc0",-- -580
x"fba60",-- -1114
x"01900",-- 400
x"01fd0",-- 509
x"fdc70",-- -569
x"02640",-- 612
x"04e00",-- 1248
x"022f0",-- 559
x"06080",-- 1544
x"051c0",-- 1308
x"07630",-- 1891
x"09ea0",-- 2538
x"09100",-- 2320
x"0c4a0",-- 3146
x"0dfd0",-- 3581
x"0c5f0",-- 3167
x"097e0",-- 2430
x"0f060",-- 3846
x"13600",-- 4960
x"0dec0",-- 3564
x"0bc90",-- 3017
x"15870",-- 5511
x"17e10",-- 6113
x"0b900",-- 2960
x"0cfc0",-- 3324
x"18c80",-- 6344
x"11a80",-- 4520
x"0cd60",-- 3286
x"14ff0",-- 5375
x"167f0",-- 5759
x"12b30",-- 4787
x"10520",-- 4178
x"13420",-- 4930
x"150e0",-- 5390
x"11da0",-- 4570
x"0eff0",-- 3839
x"0f6d0",-- 3949
x"10a20",-- 4258
x"0c630",-- 3171
x"07150",-- 1813
x"094a0",-- 2378
x"08280",-- 2088
x"016c0",-- 364
x"00ef0",-- 239
x"03590",-- 857
x"fee90",-- -279
x"f7160",-- -2282
x"f58b0",-- -2677
x"f6f30",-- -2317
x"f1ea0",-- -3606
x"ec5a0",-- -5030
x"eee80",-- -4376
x"efbd0",-- -4163
x"ea560",-- -5546
x"e8b00",-- -5968
x"eb7c0",-- -5252
x"eb470",-- -5305
x"e7dd0",-- -6179
x"ea740",-- -5516
x"efb00",-- -4176
x"f03f0",-- -4033
x"ef160",-- -4330
x"f1ed0",-- -3603
x"f5e70",-- -2585
x"f4e90",-- -2839
x"f6440",-- -2492
x"fad50",-- -1323
x"fcb10",-- -847
x"fb9e0",-- -1122
x"fc1b0",-- -997
x"fe2d0",-- -467
x"fe070",-- -505
x"fd270",-- -729
x"fd4e0",-- -690
x"fe490",-- -439
x"fe690",-- -407
x"fc3f0",-- -961
x"fbbd0",-- -1091
x"fb480",-- -1208
x"f8340",-- -1996
x"f6d20",-- -2350
x"f6690",-- -2455
x"f6320",-- -2510
x"f5dd0",-- -2595
x"f4d50",-- -2859
x"f3a90",-- -3159
x"f31a0",-- -3302
x"f2890",-- -3447
x"f3890",-- -3191
x"f6c10",-- -2367
x"f8a70",-- -1881
x"f83c0",-- -1988
x"f9830",-- -1661
x"fb560",-- -1194
x"fbd60",-- -1066
x"ff220",-- -222
x"011c0",-- 284
x"02520",-- 594
x"048c0",-- 1164
x"052b0",-- 1323
x"09ea0",-- 2538
x"0a550",-- 2645
x"048a0",-- 1162
x"08e80",-- 2280
x"10c00",-- 4288
x"09b80",-- 2488
x"09240",-- 2340
x"13510",-- 4945
x"0d090",-- 3337
x"07220",-- 1826
x"0db00",-- 3504
x"10cc0",-- 4300
x"0af90",-- 2809
x"095b0",-- 2395
x"0e6b0",-- 3691
x"0eaa0",-- 3754
x"0b130",-- 2835
x"06340",-- 1588
x"0bbc0",-- 3004
x"11590",-- 4441
x"0be40",-- 3044
x"0a390",-- 2617
x"11b90",-- 4537
x"12220",-- 4642
x"0d1c0",-- 3356
x"0e8c0",-- 3724
x"11bf0",-- 4543
x"14720",-- 5234
x"11ce0",-- 4558
x"12280",-- 4648
x"165f0",-- 5727
x"12610",-- 4705
x"0c700",-- 3184
x"0c180",-- 3096
x"0ceb0",-- 3307
x"0a720",-- 2674
x"07e70",-- 2023
x"08730",-- 2163
x"05a80",-- 1448
x"00620",-- 98
x"fd760",-- -650
x"fcda0",-- -806
x"f85a0",-- -1958
x"f13e0",-- -3778
x"f0440",-- -4028
x"f2230",-- -3549
x"ee440",-- -4540
x"e9c00",-- -5696
x"ea300",-- -5584
x"e85a0",-- -6054
x"e56f0",-- -6801
x"e6830",-- -6525
x"eae80",-- -5400
x"ebd40",-- -5164
x"eaee0",-- -5394
x"ed0c0",-- -4852
x"f1220",-- -3806
x"f2a70",-- -3417
x"f2a70",-- -3417
x"f6480",-- -2488
x"f9950",-- -1643
x"fa990",-- -1383
x"fc6c0",-- -916
x"ffc20",-- -62
x"00980",-- 152
x"ffc70",-- -57
x"00640",-- 100
x"01900",-- 400
x"01990",-- 409
x"00800",-- 128
x"00800",-- 128
x"00910",-- 145
x"fe9b0",-- -357
x"fb7b0",-- -1157
x"fa7b0",-- -1413
x"f9ae0",-- -1618
x"f74a0",-- -2230
x"f6610",-- -2463
x"f6e10",-- -2335
x"f6530",-- -2477
x"f40c0",-- -3060
x"f2930",-- -3437
x"f3560",-- -3242
x"f41e0",-- -3042
x"f3040",-- -3324
x"f2ca0",-- -3382
x"f54d0",-- -2739
x"f7e00",-- -2080
x"f9d00",-- -1584
x"fafc0",-- -1284
x"fbbd0",-- -1091
x"fcb10",-- -847
x"feed0",-- -275
x"018a0",-- 394
x"036f0",-- 879
x"03a40",-- 932
x"048c0",-- 1164
x"06550",-- 1621
x"07830",-- 1923
x"08e50",-- 2277
x"09bc0",-- 2492
x"09c10",-- 2497
x"071d0",-- 1821
x"07380",-- 1848
x"0d9c0",-- 3484
x"0e540",-- 3668
x"03da0",-- 986
x"07b50",-- 1973
x"111f0",-- 4383
x"086d0",-- 2157
x"03100",-- 784
x"0c2d0",-- 3117
x"10190",-- 4121
x"06430",-- 1603
x"03650",-- 869
x"10040",-- 4100
x"0efc0",-- 3836
x"04440",-- 1092
x"094f0",-- 2383
x"13be0",-- 5054
x"0f420",-- 3906
x"09b00",-- 2480
x"11c90",-- 4553
x"13830",-- 4995
x"0ef70",-- 3831
x"11330",-- 4403
x"12590",-- 4697
x"11590",-- 4441
x"10f90",-- 4345
x"0d310",-- 3377
x"09c20",-- 2498
x"0b580",-- 2904
x"0bb80",-- 3000
x"08630",-- 2147
x"078d0",-- 1933
x"07a30",-- 1955
x"035b0",-- 859
x"fe7d0",-- -387
x"feb40",-- -332
x"fcb90",-- -839
x"f5d60",-- -2602
x"f3b10",-- -3151
x"f6620",-- -2462
x"f2fc0",-- -3332
x"ede80",-- -4632
x"ef930",-- -4205
x"eef30",-- -4365
x"e9a20",-- -5726
x"e9330",-- -5837
x"ee290",-- -4567
x"eed00",-- -4400
x"ed270",-- -4825
x"ef2e0",-- -4306
x"f2f80",-- -3336
x"f3150",-- -3307
x"f1fb0",-- -3589
x"f5a40",-- -2652
x"f8570",-- -1961
x"f8320",-- -1998
x"f9e00",-- -1568
x"fe690",-- -407
x"ff540",-- -172
x"fdf90",-- -519
x"ff360",-- -202
x"00a00",-- 160
x"00460",-- 70
x"ff070",-- -249
x"00580",-- 88
x"00f90",-- 249
x"ff800",-- -128
x"fd8d0",-- -627
x"fc1b0",-- -997
x"faa00",-- -1376
x"f8a50",-- -1883
x"f9480",-- -1720
x"fa160",-- -1514
x"f9330",-- -1741
x"f7400",-- -2240
x"f6190",-- -2535
x"f6320",-- -2510
x"f6d20",-- -2350
x"f6980",-- -2408
x"f75c0",-- -2212
x"f94a0",-- -1718
x"f94d0",-- -1715
x"fa3a0",-- -1478
x"fc390",-- -967
x"fb880",-- -1144
x"fb510",-- -1199
x"fd590",-- -679
x"00480",-- 72
x"02ff0",-- 767
x"03880",-- 904
x"02910",-- 657
x"031d0",-- 797
x"04bb0",-- 1211
x"03900",-- 912
x"03b50",-- 949
x"04d10",-- 1233
x"05670",-- 1383
x"076a0",-- 1898
x"05450",-- 1349
x"03a30",-- 931
x"062a0",-- 1578
x"06f70",-- 1783
x"03010",-- 769
x"018a0",-- 394
x"08080",-- 2056
x"08d70",-- 2263
x"02260",-- 550
x"043a0",-- 1082
x"07e40",-- 2020
x"05c90",-- 1481
x"04110",-- 1041
x"06c70",-- 1735
x"08aa0",-- 2218
x"05f80",-- 1528
x"067b0",-- 1659
x"08f70",-- 2295
x"08660",-- 2150
x"06dc0",-- 1756
x"07bc0",-- 1980
x"0aac0",-- 2732
x"08d10",-- 2257
x"08e30",-- 2275
x"0ca00",-- 3232
x"0abe0",-- 2750
x"08840",-- 2180
x"0b590",-- 2905
x"0c7f0",-- 3199
x"09170",-- 2327
x"084b0",-- 2123
x"09c40",-- 2500
x"0a820",-- 2690
x"0a5f0",-- 2655
x"0a590",-- 2649
x"0a690",-- 2665
x"08be0",-- 2238
x"067a0",-- 1658
x"05760",-- 1398
x"03f40",-- 1012
x"02200",-- 544
x"00dc0",-- 220
x"ff8b0",-- -117
x"fdb50",-- -587
x"fc530",-- -941
x"fb770",-- -1161
x"f9c90",-- -1591
x"f7e40",-- -2076
x"f6be0",-- -2370
x"f6570",-- -2473
x"f6160",-- -2538
x"f63c0",-- -2500
x"f6530",-- -2477
x"f60f0",-- -2545
x"f5700",-- -2704
x"f54a0",-- -2742
x"f62b0",-- -2517
x"f6ca0",-- -2358
x"f73b0",-- -2245
x"f87d0",-- -1923
x"f9590",-- -1703
x"f94f0",-- -1713
x"fa140",-- -1516
x"fa5d0",-- -1443
x"f9cb0",-- -1589
x"f92f0",-- -1745
x"f8b90",-- -1863
x"f9420",-- -1726
x"f8fc0",-- -1796
x"f88f0",-- -1905
x"f89e0",-- -1890
x"f8760",-- -1930
x"f8390",-- -1991
x"f82d0",-- -2003
x"f9310",-- -1743
x"f8cf0",-- -1841
x"f90e0",-- -1778
x"f9950",-- -1643
x"f9d80",-- -1576
x"fa670",-- -1433
x"facf0",-- -1329
x"faeb0",-- -1301
x"fa8a0",-- -1398
x"fc2d0",-- -979
x"fddf0",-- -545
x"fee10",-- -287
x"fef00",-- -272
x"fe7d0",-- -387
x"fefa0",-- -262
x"ff440",-- -188
x"ff7c0",-- -132
x"ffdf0",-- -33
x"00370",-- 55
x"ffa60",-- -90
x"ffab0",-- -85
x"00ad0",-- 173
x"012b0",-- 299
x"00e80",-- 232
x"006e0",-- 110
x"015d0",-- 349
x"01f90",-- 505
x"02030",-- 515
x"02b40",-- 692
x"03b30",-- 947
x"03a40",-- 932
x"03360",-- 822
x"04030",-- 1027
x"04de0",-- 1246
x"047f0",-- 1151
x"045d0",-- 1117
x"04f00",-- 1264
x"05100",-- 1296
x"04a90",-- 1193
x"05130",-- 1299
x"05400",-- 1344
x"05060",-- 1286
x"04d40",-- 1236
x"04990",-- 1177
x"04940",-- 1172
x"04490",-- 1097
x"047a0",-- 1146
x"04170",-- 1047
x"04000",-- 1024
x"04370",-- 1079
x"03f60",-- 1014
x"04070",-- 1031
x"043f0",-- 1087
x"04980",-- 1176
x"04750",-- 1141
x"04e50",-- 1253
x"058f0",-- 1423
x"060a0",-- 1546
x"06700",-- 1648
x"06ed0",-- 1773
x"07b20",-- 1970
x"07e00",-- 2016
x"08840",-- 2180
x"09790",-- 2425
x"09ee0",-- 2542
x"09cc0",-- 2508
x"09d30",-- 2515
x"09c40",-- 2500
x"09270",-- 2343
x"085c0",-- 2140
x"07e70",-- 2023
x"074a0",-- 1866
x"06050",-- 1541
x"04f90",-- 1273
x"04210",-- 1057
x"02fc0",-- 764
x"01ae0",-- 430
x"00320",-- 50
x"ff3d0",-- -195
x"fe0d0",-- -499
x"fd240",-- -732
x"fc910",-- -879
x"fc0f0",-- -1009
x"fb740",-- -1164
x"fa850",-- -1403
x"fa440",-- -1468
x"f9e20",-- -1566
x"f8e40",-- -1820
x"f84e0",-- -1970
x"f82b0",-- -2005
x"f78d0",-- -2163
x"f7330",-- -2253
x"f6da0",-- -2342
x"f6cd0",-- -2355
x"f6580",-- -2472
x"f59a0",-- -2662
x"f54f0",-- -2737
x"f54d0",-- -2739
x"f51f0",-- -2785
x"f4c60",-- -2874
x"f4f20",-- -2830
x"f5750",-- -2699
x"f5680",-- -2712
x"f5520",-- -2734
x"f5bd0",-- -2627
x"f65c0",-- -2468
x"f6b60",-- -2378
x"f7160",-- -2282
x"f8190",-- -2023
x"f8cb0",-- -1845
x"f9340",-- -1740
x"f9f80",-- -1544
x"fb150",-- -1259
x"fba60",-- -1114
x"fc390",-- -967
x"fd2c0",-- -724
x"fdab0",-- -597
x"fe3e0",-- -450
x"fed50",-- -299
x"ff760",-- -138
x"fff10",-- -15
x"003f0",-- 63
x"00a80",-- 168
x"00f70",-- 247
x"018d0",-- 397
x"02070",-- 519
x"02610",-- 609
x"02c50",-- 709
x"031f0",-- 799
x"03b20",-- 946
x"040c0",-- 1036
x"04730",-- 1139
x"04d90",-- 1241
x"05260",-- 1318
x"058f0",-- 1423
x"05fb0",-- 1531
x"063e0",-- 1598
x"063c0",-- 1596
x"06ae0",-- 1710
x"06d10",-- 1745
x"06be0",-- 1726
x"06c20",-- 1730
x"06bb0",-- 1723
x"06640",-- 1636
x"05e40",-- 1508
x"05d60",-- 1494
x"05b80",-- 1464
x"05580",-- 1368
x"04d10",-- 1233
x"04ca0",-- 1226
x"04980",-- 1176
x"04170",-- 1047
x"03f40",-- 1012
x"04230",-- 1059
x"03f80",-- 1016
x"03da0",-- 986
x"04080",-- 1032
x"04070",-- 1031
x"042a0",-- 1066
x"042a0",-- 1066
x"049d0",-- 1181
x"05080",-- 1288
x"056f0",-- 1391
x"05b20",-- 1458
x"05fe0",-- 1534
x"06b60",-- 1718
x"073f0",-- 1855
x"07860",-- 1926
x"079f0",-- 1951
x"078a0",-- 1930
x"07030",-- 1795
x"06370",-- 1591
x"05c70",-- 1479
x"05470",-- 1351
x"04370",-- 1079
x"03100",-- 784
x"02280",-- 552
x"012e0",-- 302
x"ffe50",-- -27
x"feeb0",-- -277
x"fdee0",-- -530
x"fd160",-- -746
x"fc250",-- -987
x"fb920",-- -1134
x"fba10",-- -1119
x"fb2a0",-- -1238
x"fad90",-- -1319
x"fa9b0",-- -1381
x"fa960",-- -1386
x"fa200",-- -1504
x"f9fd0",-- -1539
x"f9ef0",-- -1553
x"f9970",-- -1641
x"f9900",-- -1648
x"f93e0",-- -1730
x"f9740",-- -1676
x"f93e0",-- -1730
x"f8be0",-- -1858
x"f8670",-- -1945
x"f82d0",-- -2003
x"f7f90",-- -2055
x"f7830",-- -2173
x"f7a80",-- -2136
x"f7dd0",-- -2083
x"f7810",-- -2175
x"f7a10",-- -2143
x"f7e70",-- -2073
x"f7fb0",-- -2053
x"f82a0",-- -2006
x"f8850",-- -1915
x"f9150",-- -1771
x"f9970",-- -1641
x"fa140",-- -1516
x"fac00",-- -1344
x"fb680",-- -1176
x"fbb70",-- -1097
x"fc230",-- -989
x"fcfd0",-- -771
x"fd900",-- -624
x"fdfd0",-- -515
x"fe8c0",-- -372
x"ff470",-- -185
x"ffb20",-- -78
x"00050",-- 5
x"00ad0",-- 173
x"010e0",-- 270
x"01590",-- 345
x"01bd0",-- 445
x"02390",-- 569
x"02b60",-- 694
x"02d70",-- 727
x"031d0",-- 797
x"03620",-- 866
x"037c0",-- 892
x"038d0",-- 909
x"03b80",-- 952
x"04190",-- 1049
x"03ee0",-- 1006
x"03f80",-- 1016
x"04300",-- 1072
x"04120",-- 1042
x"04000",-- 1024
x"03dd0",-- 989
x"03da0",-- 986
x"038f0",-- 911
x"03450",-- 837
x"03440",-- 836
x"03270",-- 807
x"02f00",-- 752
x"027d0",-- 637
x"02670",-- 615
x"022b0",-- 555
x"01ba0",-- 442
x"01830",-- 387
x"01630",-- 355
x"01420",-- 322
x"00e80",-- 232
x"00c50",-- 197
x"00ac0",-- 172
x"00960",-- 150
x"00440",-- 68
x"00200",-- 32
x"006c0",-- 108
x"00620",-- 98
x"00730",-- 115
x"00c30",-- 195
x"01090",-- 265
x"01180",-- 280
x"014e0",-- 334
x"01a40",-- 420
x"01e20",-- 482
x"02140",-- 532
x"02410",-- 577
x"02e50",-- 741
x"03630",-- 867
x"03ab0",-- 939
x"03e70",-- 999
x"04660",-- 1126
x"04cd0",-- 1229
x"052b0",-- 1323
x"05c10",-- 1473
x"05ce0",-- 1486
x"05e90",-- 1513
x"058a0",-- 1418
x"051d0",-- 1309
x"04ef0",-- 1263
x"04690",-- 1129
x"03f30",-- 1011
x"03420",-- 834
x"02c30",-- 707
x"01ef0",-- 495
x"01290",-- 297
x"006e0",-- 110
x"ff9c0",-- -100
x"fee30",-- -285
x"fe3a0",-- -454
x"fe070",-- -505
x"fdd60",-- -554
x"fd860",-- -634
x"fd4f0",-- -689
x"fd530",-- -685
x"fcda0",-- -806
x"fc870",-- -889
x"fc8e0",-- -882
x"fc690",-- -919
x"fc300",-- -976
x"fc110",-- -1007
x"fbf40",-- -1036
x"fbe20",-- -1054
x"fbc90",-- -1079
x"fb5e0",-- -1186
x"fb010",-- -1279
x"fac10",-- -1343
x"fa750",-- -1419
x"fa2b0",-- -1493
x"fa2b0",-- -1493
x"fa0a0",-- -1526
x"f9bc0",-- -1604
x"f9850",-- -1659
x"f9830",-- -1661
x"f96d0",-- -1683
x"f98d0",-- -1651
x"f9a60",-- -1626
x"f9f10",-- -1551
x"fa460",-- -1466
x"fa8e0",-- -1394
x"fb110",-- -1263
x"fb570",-- -1193
x"fbd00",-- -1072
x"fc160",-- -1002
x"fcc10",-- -831
x"fd6f0",-- -657
x"fdf10",-- -527
x"fe9b0",-- -357
x"ff1d0",-- -227
x"ffb80",-- -72
x"00210",-- 33
x"00cb0",-- 203
x"014f0",-- 335
x"01c60",-- 454
x"023e0",-- 574
x"029d0",-- 669
x"03100",-- 784
x"03770",-- 887
x"03c60",-- 966
x"03fd0",-- 1021
x"042a0",-- 1066
x"044d0",-- 1101
x"046c0",-- 1132
x"048a0",-- 1162
x"04910",-- 1169
x"047b0",-- 1147
x"046e0",-- 1134
x"043f0",-- 1087
x"03fd0",-- 1021
x"03c10",-- 961
x"03880",-- 904
x"03330",-- 819
x"02d20",-- 722
x"028e0",-- 654
x"023f0",-- 575
x"01f30",-- 499
x"01b50",-- 437
x"01600",-- 352
x"01090",-- 265
x"00d90",-- 217
x"008c0",-- 140
x"005d0",-- 93
x"00370",-- 55
x"00000",-- 0
x"ffc90",-- -55
x"ff950",-- -107
x"ff590",-- -167
x"ff1f0",-- -225
x"fefa0",-- -262
x"febb0",-- -325
x"fe8c0",-- -372
x"fe760",-- -394
x"fe4d0",-- -435
x"fe1e0",-- -482
x"fe050",-- -507
x"fe000",-- -512
x"fde40",-- -540
x"fdf60",-- -522
x"fe170",-- -489
x"fe430",-- -445
x"fe700",-- -400
x"fe850",-- -379
x"fef80",-- -264
x"ff330",-- -205
x"ff670",-- -153
x"ffd50",-- -43
x"00480",-- 72
x"00a20",-- 162
x"00fc0",-- 252
x"01740",-- 372
x"01ec0",-- 492
x"025f0",-- 607
x"02d20",-- 722
x"03450",-- 837
x"03ce0",-- 974
x"042b0",-- 1067
x"04890",-- 1161
x"05040",-- 1284
x"05440",-- 1348
x"05600",-- 1376
x"05600",-- 1376
x"05560",-- 1366
x"051c0",-- 1308
x"04dc0",-- 1244
x"048c0",-- 1164
x"04320",-- 1074
x"03b30",-- 947
x"03210",-- 801
x"02a00",-- 672
x"02050",-- 517
x"01670",-- 359
x"00d20",-- 210
x"00670",-- 103
x"ffdb0",-- -37
x"ff860",-- -122
x"ff380",-- -200
x"fefd0",-- -259
x"febb0",-- -325
x"fe660",-- -410
x"fe2b0",-- -469
x"fdea0",-- -534
x"fdb80",-- -584
x"fd6a0",-- -662
x"fd530",-- -685
x"fd020",-- -766
x"fca20",-- -862
x"fc710",-- -911
x"fc300",-- -976
x"fbd30",-- -1069
x"fb940",-- -1132
x"fb540",-- -1196
x"fb020",-- -1278
x"fae60",-- -1306
x"fac60",-- -1338
x"fab40",-- -1356
x"faa30",-- -1373
x"faa50",-- -1371
x"faa30",-- -1373
x"faca0",-- -1334
x"fb1a0",-- -1254
x"fb4d0",-- -1203
x"fb9c0",-- -1124
x"fc050",-- -1019
x"fc760",-- -906
x"fcda0",-- -806
x"fd440",-- -700
x"fdbf0",-- -577
x"fe140",-- -492
x"fe8a0",-- -374
x"ff010",-- -255
x"ff580",-- -168
x"ffce0",-- -50
x"00110",-- 17
x"00670",-- 103
x"00a70",-- 167
x"00ef0",-- 239
x"01290",-- 297
x"01630",-- 355
x"01970",-- 407
x"01bf0",-- 447
x"02070",-- 519
x"02160",-- 534
x"023c0",-- 572
x"023c0",-- 572
x"024e0",-- 590
x"02340",-- 564
x"02320",-- 562
x"024b0",-- 587
x"02350",-- 565
x"02460",-- 582
x"022a0",-- 554
x"02250",-- 549
x"020f0",-- 527
x"01f90",-- 505
x"01f60",-- 502
x"01e90",-- 489
x"01db0",-- 475
x"01b70",-- 439
x"019f0",-- 415
x"019e0",-- 414
x"016a0",-- 362
x"01420",-- 322
x"01290",-- 297
x"00f90",-- 249
x"00e30",-- 227
x"00a50",-- 165
x"00800",-- 128
x"005a0",-- 90
x"00280",-- 40
x"00070",-- 7
x"fff80",-- -8
x"fff90",-- -7
x"ffc60",-- -58
x"ffb50",-- -75
x"ffc20",-- -62
x"ffcc0",-- -52
x"ffbf0",-- -65
x"ffd60",-- -42
x"fff30",-- -13
x"fffb0",-- -5
x"000f0",-- 15
x"00280",-- 40
x"005a0",-- 90
x"007b0",-- 123
x"00960",-- 150
x"00dc0",-- 220
x"01100",-- 272
x"013b0",-- 315
x"01860",-- 390
x"01ec0",-- 492
x"02260",-- 550
x"02580",-- 600
x"02d20",-- 722
x"031a0",-- 794
x"03590",-- 857
x"039a0",-- 922
x"03b00",-- 944
x"03c10",-- 961
x"03a60",-- 934
x"03920",-- 914
x"036f0",-- 879
x"03350",-- 821
x"02de0",-- 734
x"02870",-- 647
x"024d0",-- 589
x"01ae0",-- 430
x"01420",-- 322
x"00d70",-- 215
x"006b0",-- 107
x"fff40",-- -12
x"ff8b0",-- -117
x"ff6a0",-- -150
x"ff1d0",-- -227
x"fee40",-- -284
x"fe8c0",-- -372
x"fe6b0",-- -405
x"fe480",-- -440
x"fdf30",-- -525
x"fdd30",-- -557
x"fdbc0",-- -580
x"fd8b0",-- -629
x"fd560",-- -682
x"fd3d0",-- -707
x"fd160",-- -746
x"fcf70",-- -777
x"fcb40",-- -844
x"fc8f0",-- -881
x"fc8a0",-- -886
x"fc4d0",-- -947
x"fc340",-- -972
x"fc260",-- -986
x"fc1c0",-- -996
x"fbfd0",-- -1027
x"fc020",-- -1022
x"fc1c0",-- -996
x"fc1c0",-- -996
x"fc3f0",-- -961
x"fc5a0",-- -934
x"fc9b0",-- -869
x"fcc80",-- -824
x"fcf00",-- -784
x"fd4e0",-- -690
x"fd810",-- -639
x"fdb20",-- -590
x"fdf40",-- -524
x"fe520",-- -430
x"fe7f0",-- -385
x"feb60",-- -330
x"ff040",-- -252
x"ff310",-- -207
x"ff5d0",-- -163
x"ff970",-- -105
x"ffce0",-- -50
x"000c0",-- 12
x"002f0",-- 47
x"00520",-- 82
x"00aa0",-- 170
x"00e60",-- 230
x"00fc0",-- 252
x"01350",-- 309
x"01800",-- 384
x"018a0",-- 394
x"01ab0",-- 427
x"01db0",-- 475
x"01ee0",-- 494
x"01fb0",-- 507
x"020a0",-- 522
x"020a0",-- 522
x"02020",-- 514
x"02000",-- 512
x"01ec0",-- 492
x"01e20",-- 482
x"01ec0",-- 492
x"01df0",-- 479
x"01c40",-- 452
x"01c40",-- 452
x"01a40",-- 420
x"019c0",-- 412
x"01900",-- 400
x"01760",-- 374
x"01620",-- 354
x"01580",-- 344
x"01510",-- 337
x"011c0",-- 284
x"011a0",-- 282
x"00f40",-- 244
x"00e80",-- 232
x"00d40",-- 212
x"00bc0",-- 188
x"00bc0",-- 188
x"00910",-- 145
x"00910",-- 145
x"00800",-- 128
x"007f0",-- 127
x"00640",-- 100
x"004d0",-- 77
x"005d0",-- 93
x"005d0",-- 93
x"005d0",-- 93
x"00670",-- 103
x"008e0",-- 142
x"009d0",-- 157
x"00a00",-- 160
x"00ca0",-- 202
x"00ef0",-- 239
x"01210",-- 289
x"01450",-- 325
x"016a0",-- 362
x"01a60",-- 422
x"01d00",-- 464
x"01f60",-- 502
x"02320",-- 562
x"02730",-- 627
x"02870",-- 647
x"02a30",-- 675
x"02d90",-- 729
x"02e00",-- 736
x"02d70",-- 727
x"02d10",-- 721
x"02b90",-- 697
x"02850",-- 645
x"02550",-- 597
x"02140",-- 532
x"01cb0",-- 459
x"01850",-- 389
x"01240",-- 292
x"00c80",-- 200
x"00780",-- 120
x"00000",-- 0
x"ffa40",-- -92
x"ff6f0",-- -145
x"ff170",-- -233
x"feb20",-- -334
x"fe8a0",-- -374
x"fe5d0",-- -419
x"fe0a0",-- -502
x"fddf0",-- -545
x"fdb50",-- -587
x"fd770",-- -649
x"fd3d0",-- -707
x"fd1f0",-- -737
x"fd060",-- -762
x"fced0",-- -787
x"fca70",-- -857
x"fc910",-- -879
x"fc8a0",-- -886
x"fc660",-- -922
x"fc430",-- -957
x"fc350",-- -971
x"fc2a0",-- -982
x"fc160",-- -1002
x"fc1e0",-- -994
x"fc260",-- -986
x"fc440",-- -956
x"fc5c0",-- -932
x"fc670",-- -921
x"fc9e0",-- -866
x"fce30",-- -797
x"fd040",-- -764
x"fd450",-- -699
x"fd9a0",-- -614
x"fde00",-- -544
x"fe1b0",-- -485
x"fe690",-- -407
x"fec00",-- -320
x"ff090",-- -247
x"ff450",-- -187
x"ffa60",-- -90
x"00020",-- 2
x"00480",-- 72
x"008f0",-- 143
x"00d90",-- 217
x"01170",-- 279
x"01420",-- 322
x"018d0",-- 397
x"01ba0",-- 442
x"01f90",-- 505
x"021c0",-- 540
x"023a0",-- 570
x"02670",-- 615
x"027f0",-- 639
x"02890",-- 649
x"029d0",-- 669
x"02cc0",-- 716
x"02b20",-- 690
x"02ca0",-- 714
x"02d40",-- 724
x"02b60",-- 694
x"029e0",-- 670
x"02940",-- 660
x"02820",-- 642
x"025c0",-- 604
x"02530",-- 595
x"022d0",-- 557
x"02120",-- 530
x"01ec0",-- 492
x"01c20",-- 450
x"019c0",-- 412
x"01760",-- 374
x"014a0",-- 330
x"01150",-- 277
x"00fa0",-- 250
x"00d20",-- 210
x"00a50",-- 165
x"00840",-- 132
x"004b0",-- 75
x"002b0",-- 43
x"00020",-- 2
x"ffe50",-- -27
x"ffbc0",-- -68
x"ffa30",-- -93
x"ff940",-- -108
x"ff740",-- -140
x"ff790",-- -135
x"ff530",-- -173
x"ff510",-- -175
x"ff3f0",-- -193
x"ff350",-- -203
x"ff450",-- -187
x"ff440",-- -188
x"ff4f0",-- -177
x"ff4e0",-- -178
x"ff650",-- -155
x"ff6f0",-- -145
x"ff7c0",-- -132
x"ff7e0",-- -130
x"ffa10",-- -95
x"ffc20",-- -62
x"ffc90",-- -55
x"ffdd0",-- -35
x"fff10",-- -15
x"00070",-- 7
x"00000",-- 0
x"00210",-- 33
x"002b0",-- 43
x"002a0",-- 42
x"002f0",-- 47
x"00440",-- 68
x"00520",-- 82
x"00460",-- 70
x"00410",-- 65
x"004e0",-- 78
x"003a0",-- 58
x"002b0",-- 43
x"00320",-- 50
x"001e0",-- 30
x"00190",-- 25
x"00000",-- 0
x"ffea0",-- -22
x"ffe40",-- -28
x"ffd50",-- -43
x"ffb20",-- -78
x"ff970",-- -105
x"ff940",-- -108
x"ff810",-- -127
x"ff530",-- -173
x"ff540",-- -172
x"ff4e0",-- -178
x"ff310",-- -207
x"ff1d0",-- -227
x"ff170",-- -233
x"ff180",-- -232
x"fefd0",-- -259
x"fef70",-- -265
x"feeb0",-- -277
x"fee30",-- -285
x"fecb0",-- -309
x"fec50",-- -315
x"fecf0",-- -305
x"fecb0",-- -309
x"feb90",-- -327
x"febe0",-- -322
x"fee40",-- -284
x"fed20",-- -302
x"fede0",-- -290
x"ff040",-- -252
x"ff040",-- -252
x"ff150",-- -235
x"ff1c0",-- -228
x"ff470",-- -185
x"ff5d0",-- -163
x"ff5d0",-- -163
x"ff810",-- -127
x"ff950",-- -107
x"ffad0",-- -83
x"ffad0",-- -83
x"ffe50",-- -27
x"00020",-- 2
x"00120",-- 18
x"00340",-- 52
x"00530",-- 83
x"00800",-- 128
x"007a0",-- 122
x"00960",-- 150
x"00ac0",-- 172
x"00c80",-- 200
x"00cf0",-- 207
x"00e40",-- 228
x"00ff0",-- 255
x"00ff0",-- 255
x"010e0",-- 270
x"01130",-- 275
x"01270",-- 295
x"011f0",-- 287
x"011a0",-- 282
x"01100",-- 272
x"01180",-- 280
x"01090",-- 265
x"00f50",-- 245
x"01030",-- 259
x"00f90",-- 249
x"00ef0",-- 239
x"00e10",-- 225
x"00d50",-- 213
x"00bc0",-- 188
x"00b60",-- 182
x"00ac0",-- 172
x"008f0",-- 143
x"00760",-- 118
x"005f0",-- 95
x"00520",-- 82
x"004b0",-- 75
x"00350",-- 53
x"00120",-- 18
x"00000",-- 0
x"ffea0",-- -22
x"ffce0",-- -50
x"ffc90",-- -55
x"ffa10",-- -95
x"ff8a0",-- -118
x"ff7c0",-- -132
x"ff770",-- -137
x"ff6c0",-- -148
x"ff580",-- -168
x"ff580",-- -168
x"ff470",-- -185
x"ff4a0",-- -182
x"ff310",-- -207
x"ff300",-- -208
x"ff440",-- -188
x"ff2e0",-- -210
x"ff240",-- -220
x"ff310",-- -207
x"ff2e0",-- -210
x"ff350",-- -203
x"ff440",-- -188
x"ff510",-- -175
x"ff540",-- -172
x"ff670",-- -153
x"ff850",-- -123
x"ff800",-- -128
x"ff8a0",-- -118
x"ff900",-- -112
x"ffa40",-- -92
x"ffb50",-- -75
x"ffbf0",-- -65
x"ffc90",-- -55
x"ffe70",-- -25
x"ffea0",-- -22
x"ffe90",-- -23
x"00020",-- 2
x"000f0",-- 15
x"000f0",-- 15
x"001b0",-- 27
x"003a0",-- 58
x"00370",-- 55
x"003f0",-- 63
x"00520",-- 82
x"00660",-- 102
x"00640",-- 100
x"00640",-- 100
x"006b0",-- 107
x"00750",-- 117
x"00890",-- 137
x"00580",-- 88
x"00730",-- 115
x"008a0",-- 138
x"00620",-- 98
x"00730",-- 115
x"00840",-- 132
x"00760",-- 118
x"00760",-- 118
x"00840",-- 132
x"00700",-- 112
x"00710",-- 113
x"00730",-- 115
x"00700",-- 112
x"00620",-- 98
x"00570",-- 87
x"00480",-- 72
x"00440",-- 68
x"004e0",-- 78
x"00440",-- 68
x"00340",-- 52
x"00350",-- 53
x"00390",-- 57
x"00210",-- 33
x"001b0",-- 27
x"001b0",-- 27
x"00160",-- 22
x"00000",-- 0
x"00080",-- 8
x"00190",-- 25
x"000c0",-- 12
x"00050",-- 5
x"000a0",-- 10
x"00120",-- 18
x"00050",-- 5
x"00000",-- 0
x"000d0",-- 13
x"00030",-- 3
x"fff90",-- -7
x"fffb0",-- -5
x"00070",-- 7
x"fffe0",-- -2
x"fff90",-- -7
x"00080",-- 8
x"000c0",-- 12
x"fffe0",-- -2
x"00000",-- 0
x"000c0",-- 12
x"00030",-- 3
x"00000",-- 0
x"fffe0",-- -2
x"00140",-- 20
x"00050",-- 5
x"fffe0",-- -2
x"00000",-- 0
x"00000",-- 0
x"fff60",-- -10
x"ffe50",-- -27
x"fff80",-- -8
x"fff60",-- -10
x"ffea0",-- -22
x"ffe70",-- -25
x"ffdb0",-- -37
x"ffe40",-- -28
x"ffce0",-- -50
x"ffc60",-- -58
x"ffd00",-- -48
x"ffd10",-- -47
x"ffbf0",-- -65
x"ffb20",-- -78
x"ffc10",-- -63
x"ffb50",-- -75
x"ffa80",-- -88
x"ffa40",-- -92
x"ffad0",-- -83
x"ffa90",-- -87
x"ff9f0",-- -97
x"ffa30",-- -93
x"ffa90",-- -87
x"ffa30",-- -93
x"ff9f0",-- -97
x"ffa80",-- -88
x"ff9a0",-- -102
x"ffa10",-- -95
x"ff990",-- -103
x"ff990",-- -103
x"ff9c0",-- -100
x"ff950",-- -107
x"ff950",-- -107
x"ffa40",-- -92
x"ffa40",-- -92
x"ff8f0",-- -113
x"ffb30",-- -77
x"ffb00",-- -80
x"ffb30",-- -77
x"ffc70",-- -57
x"ffd10",-- -47
x"ffc90",-- -55
x"ffd10",-- -47
x"ffdf0",-- -33
x"ffdf0",-- -33
x"fff60",-- -10
x"fffd0",-- -3
x"00000",-- 0
x"00000",-- 0
x"00120",-- 18
x"00190",-- 25
x"00210",-- 33
x"00250",-- 37
x"001c0",-- 28
x"00320",-- 50
x"00410",-- 65
x"00460",-- 70
x"004e0",-- 78
x"004d0",-- 77
x"00500",-- 80
x"004e0",-- 78
x"00580",-- 88
x"005c0",-- 92
x"00670",-- 103
x"00700",-- 112
x"00670",-- 103
x"007a0",-- 122
x"006b0",-- 107
x"006c0",-- 108
x"00700",-- 112
x"00690",-- 105
x"00700",-- 112
x"00700",-- 112
x"007b0",-- 123
x"00760",-- 118
x"00710",-- 113
x"006b0",-- 107
x"00610",-- 97
x"005c0",-- 92
x"00620",-- 98
x"006e0",-- 110
x"005f0",-- 95
x"00570",-- 87
x"005a0",-- 90
x"005a0",-- 90
x"00480",-- 72
x"003c0",-- 60
x"00520",-- 82
x"00410",-- 65
x"00320",-- 50
x"00350",-- 53
x"00340",-- 52
x"00320",-- 50
x"00250",-- 37
x"001c0",-- 28
x"001b0",-- 27
x"000f0",-- 15
x"000a0",-- 10
x"000a0",-- 10
x"000d0",-- 13
x"000f0",-- 15
x"00000",-- 0
x"000a0",-- 10
x"000a0",-- 10
x"000c0",-- 12
x"00080",-- 8
x"00190",-- 25
x"00260",-- 38
x"001b0",-- 27
x"000f0",-- 15
x"000c0",-- 12
x"000d0",-- 13
x"00070",-- 7
x"000f0",-- 15
x"00190",-- 25
x"00080",-- 8
x"000d0",-- 13
x"00020",-- 2
x"00050",-- 5
x"00050",-- 5
x"fff40",-- -12
x"00020",-- 2
x"00080",-- 8
x"00070",-- 7
x"fffe0",-- -2
x"00080",-- 8
x"fffe0",-- -2
x"fff60",-- -10
x"fff80",-- -8
x"fff90",-- -7
x"00050",-- 5
x"fffe0",-- -2
x"00070",-- 7
x"00030",-- 3
x"00020",-- 2
x"00000",-- 0
x"00000",-- 0
x"00020",-- 2
x"fffd0",-- -3
x"000c0",-- 12
x"00080",-- 8
x"000f0",-- 15
x"00050",-- 5
x"00050",-- 5
x"000a0",-- 10
x"00070",-- 7
x"00000",-- 0
x"fffb0",-- -5
x"00080",-- 8
x"fffe0",-- -2
x"fff30",-- -13
x"00000",-- 0
x"fffd0",-- -3
x"fff80",-- -8
x"ffef0",-- -17
x"ffe50",-- -27
x"ffee0",-- -18
x"ffee0",-- -18
x"ffdb0",-- -37
x"ffe50",-- -27
x"ffea0",-- -22
x"ffe00",-- -32
x"ffe70",-- -25
x"ffe00",-- -32
x"ffe40",-- -28
x"ffea0",-- -22
x"fff10",-- -15
x"fff40",-- -12
x"fff80",-- -8
x"fffe0",-- -2
x"00000",-- 0
x"00000",-- 0
x"fff30",-- -13
x"fffb0",-- -5
x"00000",-- 0
x"fff40",-- -12
x"fffd0",-- -3
x"fffd0",-- -3
x"fffe0",-- -2
x"00000",-- 0
x"00000",-- 0
x"000a0",-- 10
x"000a0",-- 10
x"000a0",-- 10
x"00030",-- 3
x"000f0",-- 15
x"000f0",-- 15
x"00120",-- 18
x"00080",-- 8
x"000c0",-- 12
x"000c0",-- 12
x"000d0",-- 13
x"00190",-- 25
x"00160",-- 22
x"000d0",-- 13
x"00050",-- 5
x"000d0",-- 13
x"000d0",-- 13
x"000d0",-- 13
x"000d0",-- 13
x"000f0",-- 15
x"000a0",-- 10
x"00020",-- 2
x"00080",-- 8
x"00030",-- 3
x"00020",-- 2
x"00050",-- 5
x"00000",-- 0
x"00050",-- 5
x"00050",-- 5
x"00050",-- 5
x"00070",-- 7
x"fffe0",-- -2
x"00000",-- 0
x"00020",-- 2
x"00080",-- 8
x"00000",-- 0
x"00020",-- 2
x"00050",-- 5
x"fff80",-- -8
x"fff80",-- -8
x"fff60",-- -10
x"fff40",-- -12
x"fff10",-- -15
x"fffd0",-- -3
x"fffe0",-- -2
x"fff40",-- -12
x"fffb0",-- -5
x"fff90",-- -7
x"fff40",-- -12
x"fff80",-- -8
x"ffee0",-- -18
x"fffb0",-- -5
x"fffe0",-- -2
x"fffb0",-- -5
x"fff90",-- -7
x"fffd0",-- -3
x"00000",-- 0
x"fff40",-- -12
x"00000",-- 0
x"fffb0",-- -5
x"fffb0",-- -5
x"fffb0",-- -5
x"fff80",-- -8
x"fffd0",-- -3
x"fff80",-- -8
x"fff40",-- -12
x"fff10",-- -15
x"fff90",-- -7
x"fffe0",-- -2
x"fff40",-- -12
x"fff10",-- -15
x"fff40",-- -12
x"fff40",-- -12
x"fff80",-- -8
x"fff40",-- -12
x"fff40",-- -12
x"ffef0",-- -17
x"ffe50",-- -27
x"fff60",-- -10
x"fff80",-- -8
x"ffef0",-- -17
x"fff60",-- -10
x"00000",-- 0
x"fff80",-- -8
x"ffef0",-- -17
x"fff40",-- -12
x"fff10",-- -15
x"ffe70",-- -25
x"fff30",-- -13
x"fffe0",-- -2
x"fff10",-- -15
x"ffe70",-- -25
x"ffe40",-- -28
x"ffea0",-- -22
x"ffe50",-- -27
x"ffdb0",-- -37
x"ffda0",-- -38
x"ffd60",-- -42
x"ffd50",-- -43
x"ffd50",-- -43
x"ffda0",-- -38
x"ffe50",-- -27
x"ffe90",-- -23
x"ffdf0",-- -33
x"ffda0",-- -38
x"ffe20",-- -30
x"ffd80",-- -40
x"ffce0",-- -50
x"ffdf0",-- -33
x"ffda0",-- -38
x"ffd30",-- -45
x"ffce0",-- -50
x"ffd60",-- -42
x"ffd80",-- -40
x"ffd30",-- -45
x"ffd80",-- -40
x"ffd50",-- -43
x"ffdb0",-- -37
x"ffdb0",-- -37
x"ffe00",-- -32
x"ffda0",-- -38
x"ffd50",-- -43
x"ffd10",-- -47
x"ffe20",-- -30
x"ffe00",-- -32
x"ffdd0",-- -35
x"ffee0",-- -18
x"ffea0",-- -22
x"ffe50",-- -27
x"ffd30",-- -45
x"ffd50",-- -43
x"ffda0",-- -38
x"ffd10",-- -47
x"ffdd0",-- -35
x"ffe90",-- -23
x"ffef0",-- -17
x"ffef0",-- -17
x"fff60",-- -10
x"fff30",-- -13
x"ffef0",-- -17
x"ffee0",-- -18
x"fff80",-- -8
x"fff10",-- -15
x"fff10",-- -15
x"fff90",-- -7
x"fffb0",-- -5
x"00000",-- 0
x"00020",-- 2
x"000c0",-- 12
x"000a0",-- 10
x"00070",-- 7
x"fffd0",-- -3
x"fff80",-- -8
x"fffe0",-- -2
x"00000",-- 0
x"00080",-- 8
x"000c0",-- 12
x"00050",-- 5
x"00050",-- 5
x"00020",-- 2
x"000a0",-- 10
x"000f0",-- 15
x"000d0",-- 13
x"00110",-- 17
x"000f0",-- 15
x"00160",-- 22
x"00080",-- 8
x"000f0",-- 15
x"00000",-- 0
x"fffb0",-- -5
x"fffe0",-- -2
x"00000",-- 0
x"00080",-- 8
x"00000",-- 0
x"000c0",-- 12
x"00050",-- 5
x"00070",-- 7
x"00030",-- 3
x"00050",-- 5
x"00020",-- 2
x"00000",-- 0
x"00000",-- 0
x"00020",-- 2
x"00000",-- 0
x"fff80",-- -8
x"00000",-- 0
x"00020",-- 2
x"00020",-- 2
x"00030",-- 3
x"000d0",-- 13
x"000c0",-- 12
x"00050",-- 5
x"00070",-- 7
x"00000",-- 0
x"fffe0",-- -2
x"00000",-- 0
x"00000",-- 0
x"fffe0",-- -2
x"fffe0",-- -2
x"00000",-- 0
x"fffb0",-- -5
x"00030",-- 3
x"00050",-- 5
x"fff90",-- -7
x"fffe0",-- -2
x"fffe0",-- -2
x"fff40",-- -12
x"ffee0",-- -18
x"fff30",-- -13
x"ffea0",-- -22
x"ffe70",-- -25
x"ffe70",-- -25
x"ffe40",-- -28
x"ffec0",-- -20
x"ffea0",-- -22
x"ffe40",-- -28
x"ffea0",-- -22
x"ffea0",-- -22
x"ffdd0",-- -35
x"ffe40",-- -28
x"ffee0",-- -18
x"ffe90",-- -23
x"ffdd0",-- -35
x"ffdf0",-- -33
x"ffe00",-- -32
x"ffd50",-- -43
x"ffd50",-- -43
x"ffdb0",-- -37
x"ffe20",-- -30
x"ffe20",-- -30
x"ffe20",-- -30
x"ffdf0",-- -33
x"ffd60",-- -42
x"ffce0",-- -50
x"ffdd0",-- -35
x"ffea0",-- -22
x"ffe20",-- -30
x"ffe50",-- -27
x"ffef0",-- -17
x"ffee0",-- -18
x"ffee0",-- -18
x"ffef0",-- -17
x"fff10",-- -15
x"ffee0",-- -18
x"ffe90",-- -23
x"ffe50",-- -27
x"ffea0",-- -22
x"ffef0",-- -17
x"ffe50",-- -27
x"ffec0",-- -20
x"fffb0",-- -5
x"fff90",-- -7
x"fff30",-- -13
x"fff40",-- -12
x"fff40",-- -12
x"ffee0",-- -18
x"ffee0",-- -18
x"fff40",-- -12
x"fffb0",-- -5
x"ffea0",-- -22
x"ffee0",-- -18
x"fff60",-- -10
x"fff10",-- -15
x"fffb0",-- -5
x"00000",-- 0
x"00000",-- 0
x"00030",-- 3
x"fffe0",-- -2
x"00000",-- 0
x"fffb0",-- -5
x"fffb0",-- -5
x"fffe0",-- -2
x"00030",-- 3
x"000a0",-- 10
x"00020",-- 2
x"000a0",-- 10
x"00120",-- 18
x"00140",-- 20
x"00050",-- 5
x"000d0",-- 13
x"00110",-- 17
x"000f0",-- 15
x"00120",-- 18
x"000f0",-- 15
x"00140",-- 20
x"000a0",-- 10
x"000c0",-- 12
x"000f0",-- 15
x"00110",-- 17
x"000f0",-- 15
x"00080",-- 8
x"000c0",-- 12
x"00020",-- 2
x"000c0",-- 12
x"000c0",-- 12
x"00160",-- 22
x"00110",-- 17
x"000f0",-- 15
x"00230",-- 35
x"00190",-- 25
x"001e0",-- 30
x"00250",-- 37
x"00210",-- 33
x"00250",-- 37
x"00230",-- 35
x"00210",-- 33
x"002a0",-- 42
x"002f0",-- 47
x"00250",-- 37
x"002a0",-- 42
x"00280",-- 40
x"00260",-- 38
x"002b0",-- 43
x"001b0",-- 27
x"00280",-- 40
x"00210",-- 33
x"002b0",-- 43
x"00280",-- 40
x"00170",-- 23
x"00120",-- 18
x"000d0",-- 13
x"00080",-- 8
x"000a0",-- 10
x"00120",-- 18
x"000d0",-- 13
x"00050",-- 5
x"00000",-- 0
x"00000",-- 0
x"00020",-- 2
x"00080",-- 8
x"000c0",-- 12
x"00080",-- 8
x"00020",-- 2
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fffb0",-- -5
x"fff90",-- -7
x"00000",-- 0
x"fffb0",-- -5
x"fffd0",-- -3
x"00000",-- 0
x"fffe0",-- -2
x"fffb0",-- -5
x"fff80",-- -8
x"fffd0",-- -3
x"fffe0",-- -2
x"00000",-- 0
x"00000",-- 0
x"00020",-- 2
x"fffe0",-- -2
x"fffb0",-- -5
x"fff10",-- -15
x"fff60",-- -10
x"00000",-- 0
x"fffb0",-- -5
x"fff80",-- -8
x"fff40",-- -12
x"fff10",-- -15
x"ffef0",-- -17
x"fff40",-- -12
x"ffee0",-- -18
x"ffe70",-- -25
x"ffe70",-- -25
x"ffe50",-- -27
x"ffec0",-- -20
x"ffe20",-- -30
x"ffd80",-- -40
x"ffdf0",-- -33
x"ffe40",-- -28
x"ffe50",-- -27
x"ffe50",-- -27
x"ffea0",-- -22
x"ffec0",-- -20
x"ffe70",-- -25
x"ffdf0",-- -33
x"ffee0",-- -18
x"fff40",-- -12
x"fff40",-- -12
x"fffb0",-- -5
x"fffe0",-- -2
x"fffd0",-- -3
x"fff40",-- -12
x"fff90",-- -7
x"00000",-- 0
x"00030",-- 3
x"00030",-- 3
x"00120",-- 18
x"000f0",-- 15
x"00030",-- 3
x"00070",-- 7
x"00020",-- 2
x"00020",-- 2
x"00020",-- 2
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00050",-- 5
x"00050",-- 5
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"00080",-- 8
x"00000",-- 0
x"fffe0",-- -2
x"fffb0",-- -5
x"fff40",-- -12
x"fff90",-- -7
x"fff60",-- -10
x"00000",-- 0
x"fff90",-- -7
x"fff40",-- -12
x"fffe0",-- -2
x"fffd0",-- -3
x"fff80",-- -8
x"fffb0",-- -5
x"00000",-- 0
x"00000",-- 0
x"fff80",-- -8
x"ffea0",-- -22
x"fff30",-- -13
x"fff60",-- -10
x"fff40",-- -12
x"fff60",-- -10
x"fffb0",-- -5
x"00000",-- 0
x"00000",-- 0
x"fffd0",-- -3
x"00000",-- 0
x"00000",-- 0
x"fffe0",-- -2
x"00000",-- 0
x"00020",-- 2
x"fff80",-- -8
x"00000",-- 0
x"fff60",-- -10
x"fff10",-- -15
x"ffe50",-- -27
x"ffe50",-- -27
x"ffcc0",-- -52
x"ffd80",-- -40
x"ffa30",-- -93
x"ff940",-- -108
x"ff330",-- -205
x"fee60",-- -282
x"fe000",-- -512
x"fd530",-- -685
x"f9860",-- -1658
x"f1f20",-- -3598
x"fd670",-- -665
x"09a10",-- 2465
x"03260",-- 806
x"00670",-- 103
x"00c80",-- 200
x"01c90",-- 457
x"019c0",-- 412
x"013a0",-- 314
x"014c0",-- 332
x"ff180",-- -232
x"00a80",-- 168
x"01c90",-- 457
x"01bd0",-- 445
x"02dc0",-- 732
x"03fe0",-- 1022
x"042d0",-- 1069
x"02c50",-- 709
x"00a20",-- 162
x"00dc0",-- 220
x"010b0",-- 267
x"fe340",-- -460
x"00da0",-- 218
x"ffea0",-- -22
x"fc820",-- -894
x"ff4e0",-- -178
x"ff3f0",-- -193
x"fef80",-- -264
x"ff270",-- -217
x"fe4d0",-- -435
x"fe6c0",-- -404
x"00870",-- 135
x"00160",-- 22
x"00000",-- 0
x"01b00",-- 432
x"00520",-- 82
x"fc930",-- -877
x"ff860",-- -122
x"01ba0",-- 442
x"fda80",-- -600
x"ff0b0",-- -245
x"ffd00",-- -48
x"00850",-- 133
x"004e0",-- 78
x"fe960",-- -362
x"01a60",-- 422
x"00f50",-- 245
x"fe610",-- -415
x"00c10",-- 193
x"01a40",-- 420
x"00670",-- 103
x"00ef0",-- 239
x"01060",-- 262
x"ffbd0",-- -67
x"ff990",-- -103
x"01ce0",-- 462
x"ffc70",-- -57
x"fe850",-- -379
x"02840",-- 644
x"fee10",-- -287
x"00e40",-- 228
x"00020",-- 2
x"fd6c0",-- -660
x"017b0",-- 379
x"fe930",-- -365
x"fc0f0",-- -1009
x"00690",-- 105
x"00b10",-- 177
x"f8f50",-- -1803
x"fccd0",-- -819
x"ff1d0",-- -227
x"fb020",-- -1278
x"028e0",-- 654
x"ff710",-- -143
x"fe250",-- -475
x"04620",-- 1122
x"feb90",-- -327
x"030e0",-- 782
x"01db0",-- 475
x"fe7a0",-- -390
x"024e0",-- 590
x"04d90",-- 1241
x"01080",-- 264
x"02f40",-- 756
x"fbb20",-- -1102
x"f6c10",-- -2367
x"05e50",-- 1509
x"fd590",-- -679
x"ff630",-- -157
x"0a3c0",-- 2620
x"f5da0",-- -2598
x"02b40",-- 692
x"0ba10",-- 2977
x"f4dc0",-- -2852
x"08c80",-- 2248
x"05260",-- 1318
x"f6620",-- -2462
x"073b0",-- 1851
x"020a0",-- 522
x"fdee0",-- -530
x"01490",-- 329
x"07dd0",-- 2013
x"01710",-- 369
x"02c00",-- 704
x"0be90",-- 3049
x"f6e10",-- -2335
x"051f0",-- 1311
x"04190",-- 1049
x"f9510",-- -1711
x"07680",-- 1896
x"f7310",-- -2255
x"030d0",-- 781
x"00b20",-- 178
x"f8e10",-- -1823
x"036c0",-- 876
x"f9c70",-- -1593
x"f11a0",-- -3814
x"fd090",-- -759
x"11090",-- 4361
x"fb0e0",-- -1266
x"00a80",-- 168
x"06410",-- 1601
x"f4070",-- -3065
x"fe0c0",-- -500
x"06de0",-- 1758
x"f7160",-- -2282
x"fb420",-- -1214
x"080c0",-- 2060
x"fbec0",-- -1044
x"03d60",-- 982
x"03a10",-- 929
x"fdce0",-- -562
x"0ab10",-- 2737
x"03940",-- 916
x"f9da0",-- -1574
x"07c40",-- 1988
x"faaf0",-- -1361
x"fdb50",-- -587
x"06480",-- 1608
x"01080",-- 264
x"00d40",-- 212
x"ff580",-- -168
x"07940",-- 1940
x"f94a0",-- -1718
x"02bb0",-- 699
x"fd160",-- -746
x"f36f0",-- -3217
x"005d0",-- 93
x"f7240",-- -2268
x"00390",-- 57
x"fe550",-- -427
x"f6200",-- -2528
x"01210",-- 289
x"fda30",-- -605
x"ff5d0",-- -163
x"095e0",-- 2398
x"fe2a0",-- -470
x"066b0",-- 1643
x"07e50",-- 2021
x"f9340",-- -1740
x"01880",-- 392
x"052b0",-- 1323
x"f7980",-- -2152
x"ffbd0",-- -67
x"047d0",-- 1149
x"f7220",-- -2270
x"082f0",-- 2095
x"fac30",-- -1341
x"05e20",-- 1506
x"0d470",-- 3399
x"f5830",-- -2685
x"06890",-- 1673
x"fe080",-- -504
x"fc2a0",-- -982
x"001b0",-- 27
x"ff900",-- -112
x"fce30",-- -797
x"ff440",-- -188
x"02110",-- 529
x"fb010",-- -1279
x"0ba40",-- 2980
x"faa00",-- -1376
x"01740",-- 372
x"05060",-- 1286
x"fae90",-- -1303
x"05720",-- 1394
x"ff7e0",-- -130
x"fe170",-- -489
x"02260",-- 550
x"fbc40",-- -1084
x"fb570",-- -1193
x"05080",-- 1288
x"fe820",-- -382
x"f6390",-- -2503
x"0a8b0",-- 2699
x"01060",-- 262
x"f80f0",-- -2033
x"0c370",-- 3127
x"002f0",-- 47
x"fb240",-- -1244
x"06fc0",-- 1788
x"fee80",-- -280
x"01100",-- 272
x"046b0",-- 1131
x"fa960",-- -1386
x"039a0",-- 922
x"04a90",-- 1193
x"f7a60",-- -2138
x"023c0",-- 572
x"07380",-- 1848
x"f5f40",-- -2572
x"03b70",-- 951
x"06410",-- 1601
x"f6c60",-- -2362
x"083c0",-- 2108
x"fefa0",-- -262
x"f8480",-- -1976
x"0bd00",-- 3024
x"f9c60",-- -1594
x"fd850",-- -635
x"094f0",-- 2383
x"f84e0",-- -1970
x"01ad0",-- 429
x"011c0",-- 284
x"fe6b0",-- -405
x"018a0",-- 394
x"fcb40",-- -844
x"05100",-- 1296
x"fd450",-- -699
x"02b20",-- 690
x"fdea0",-- -534
x"ff740",-- -140
x"03380",-- 824
x"f9700",-- -1680
x"0a500",-- 2640
x"f5450",-- -2747
x"01670",-- 359
x"091f0",-- 2335
x"f0820",-- -3966
x"06370",-- 1591
x"05540",-- 1364
x"f5ec0",-- -2580
x"00340",-- 52
x"0a1b0",-- 2587
x"f99c0",-- -1636
x"fe850",-- -379
x"04e10",-- 1249
x"fe620",-- -414
x"fce40",-- -796
x"ff580",-- -168
x"045c0",-- 1116
x"fb9e0",-- -1122
x"ff920",-- -110
x"05490",-- 1353
x"fabc0",-- -1348
x"fe4d0",-- -435
x"03720",-- 882
x"fdbc0",-- -580
x"fcf30",-- -781
x"03530",-- 851
x"00d00",-- 208
x"f85d0",-- -1955
x"03240",-- 804
x"00700",-- 112
x"fad90",-- -1319
x"068c0",-- 1676
x"ffad0",-- -83
x"faf20",-- -1294
x"022f0",-- 559
x"00930",-- 147
x"01720",-- 370
x"fa5c0",-- -1444
x"ff810",-- -127
x"034a0",-- 842
x"01a60",-- 422
x"fbef0",-- -1041
x"01590",-- 345
x"01ba0",-- 442
x"f54a0",-- -2742
x"09060",-- 2310
x"027d0",-- 637
x"f8d00",-- -1840
x"043f0",-- 1087
x"00a30",-- 163
x"fcda0",-- -806
x"012b0",-- 299
x"02d70",-- 727
x"fbd00",-- -1072
x"00b60",-- 182
x"fe850",-- -379
x"ff620",-- -158
x"02940",-- 660
x"fe0a0",-- -502
x"02250",-- 549
x"002d0",-- 45
x"fa140",-- -1516
x"04dc0",-- 1244
x"ff130",-- -237
x"fdea0",-- -534
x"06370",-- 1591
x"f76f0",-- -2193
x"011f0",-- 287
x"045d0",-- 1117
x"fb250",-- -1243
x"fb2c0",-- -1236
x"06c50",-- 1733
x"fc110",-- -1007
x"fb0c0",-- -1268
x"10680",-- 4200
x"f5610",-- -2719
x"fd4e0",-- -690
x"06870",-- 1671
x"fe3c0",-- -452
x"03e90",-- 1001
x"f93b0",-- -1733
x"04350",-- 1077
x"fd1b0",-- -741
x"fc4d0",-- -947
x"ffdb0",-- -37
x"fb650",-- -1179
x"05310",-- 1329
x"00690",-- 105
x"fd010",-- -767
x"04750",-- 1141
x"ff180",-- -232
x"fe8a0",-- -374
x"022f0",-- 559
x"021c0",-- 540
x"02940",-- 660
x"fc2a0",-- -982
x"02430",-- 579
x"01740",-- 372
x"f9d10",-- -1583
x"00d70",-- 215
x"01e20",-- 482
x"02e00",-- 736
x"fbd50",-- -1067
x"fc0a0",-- -1014
x"06580",-- 1624
x"fc4b0",-- -949
x"f6910",-- -2415
x"05600",-- 1376
x"fc160",-- -1002
x"fafa0",-- -1286
x"01210",-- 289
x"febb0",-- -325
x"002f0",-- 47
x"fc0d0",-- -1011
x"06d60",-- 1750
x"007a0",-- 122
x"fd8f0",-- -625
x"04f00",-- 1264
x"007a0",-- 122
x"045f0",-- 1119
x"02d60",-- 726
x"fc300",-- -976
x"046b0",-- 1131
x"0b2e0",-- 2862
x"fb4c0",-- -1204
x"ff3f0",-- -193
x"076d0",-- 1901
x"00440",-- 68
x"f98d0",-- -1651
x"079c0",-- 1948
x"01540",-- 340
x"f47f0",-- -2945
x"0a9b0",-- 2715
x"f6ca0",-- -2358
x"08be0",-- 2238
x"fccd0",-- -819
x"ef720",-- -4238
x"154a0",-- 5450
x"edc90",-- -4663
x"026b0",-- 619
x"06b40",-- 1716
x"f4530",-- -2989
x"08ac0",-- 2220
x"fab10",-- -1359
x"054e0",-- 1358
x"00070",-- 7
x"00bc0",-- 188
x"05fd0",-- 1533
x"f31b0",-- -3301
x"12e80",-- 4840
x"00660",-- 102
x"fa550",-- -1451
x"04440",-- 1092
x"fbee0",-- -1042
x"0eca0",-- 3786
x"f1ed0",-- -3603
x"0c050",-- 3077
x"fa7d0",-- -1411
x"fd7c0",-- -644
x"12db0",-- 4827
x"e7b60",-- -6218
x"12bd0",-- 4797
x"008e0",-- 142
x"eb560",-- -5290
x"16ca0",-- 5834
x"fb650",-- -1179
x"f6850",-- -2427
x"07b00",-- 1968
x"f98f0",-- -1649
x"01350",-- 309
x"ffdf0",-- -33
x"019e0",-- 414
x"fd8f0",-- -625
x"fb950",-- -1131
x"fe3a0",-- -454
x"04660",-- 1126
x"083e0",-- 2110
x"ef020",-- -4350
x"041b0",-- 1051
x"0c180",-- 3096
x"f3a60",-- -3162
x"07ab0",-- 1963
x"05d50",-- 1493
x"f4f00",-- -2832
x"00d50",-- 213
x"09a30",-- 2467
x"fefa0",-- -262
x"f4f20",-- -2830
x"0dba0",-- 3514
x"fe490",-- -439
x"f5950",-- -2667
x"125c0",-- 4700
x"f3590",-- -3239
x"016c0",-- 364
x"05770",-- 1399
x"f1400",-- -3776
x"113d0",-- 4413
x"fe460",-- -442
x"f2730",-- -3469
x"05e20",-- 1506
x"ff4c0",-- -180
x"fd620",-- -670
x"00a20",-- 162
x"ff2c0",-- -212
x"fffb0",-- -5
x"035e0",-- 862
x"f9a90",-- -1623
x"02320",-- 562
x"03860",-- 902
x"f9b30",-- -1613
x"fdce0",-- -562
x"06910",-- 1681
x"fd800",-- -640
x"fd250",-- -731
x"02520",-- 594
x"fc200",-- -992
x"03da0",-- 986
x"fa7f0",-- -1409
x"03ba0",-- 954
x"00b90",-- 185
x"f88e0",-- -1906
x"0cff0",-- 3327
x"f71d0",-- -2275
x"ff4a0",-- -182
x"08300",-- 2096
x"f20a0",-- -3574
x"072c0",-- 1836
x"05880",-- 1416
x"f6200",-- -2528
x"03f30",-- 1011
x"00a80",-- 168
x"fc960",-- -874
x"014c0",-- 332
x"01d30",-- 467
x"fe820",-- -382
x"ff180",-- -232
x"00ad0",-- 173
x"fbad0",-- -1107
x"05c20",-- 1474
x"006e0",-- 110
x"fa110",-- -1519
x"03d50",-- 981
x"03760",-- 886
x"ffef0",-- -17
x"01290",-- 297
x"014a0",-- 330
x"faf50",-- -1291
x"06760",-- 1654
x"00e90",-- 233
x"f5830",-- -2685
x"09580",-- 2392
x"ff6d0",-- -147
x"f8d40",-- -1836
x"08410",-- 2113
x"fd240",-- -732
x"ff990",-- -103
x"030b0",-- 779
x"fd090",-- -759
x"ffd50",-- -43
x"04640",-- 1124
x"00f90",-- 249
x"fbda0",-- -1062
x"023e0",-- 574
x"ffd10",-- -47
x"ff670",-- -153
x"fff90",-- -7
x"fcf00",-- -784
x"fdcb0",-- -565
x"03b20",-- 946
x"04980",-- 1176
x"fd1a0",-- -742
x"fa800",-- -1408
x"05830",-- 1411
x"02780",-- 632
x"fb650",-- -1179
x"05a90",-- 1449
x"fe070",-- -505
x"fcad0",-- -851
x"01d00",-- 464
x"015e0",-- 350
x"02640",-- 612
x"fcff0",-- -769
x"005a0",-- 90
x"fd710",-- -655
x"01790",-- 377
x"03f90",-- 1017
x"f9270",-- -1753
x"04f20",-- 1266
x"fc5a0",-- -934
x"012e0",-- 302
x"06e60",-- 1766
x"fa490",-- -1463
x"ff090",-- -247
x"02670",-- 615
x"fd1f0",-- -737
x"07150",-- 1813
x"fc670",-- -921
x"00f70",-- 247
x"02d10",-- 721
x"f5740",-- -2700
x"0bef0",-- 3055
x"01720",-- 370
x"f75c0",-- -2212
x"03f90",-- 1017
x"021e0",-- 542
x"feac0",-- -340
x"00a70",-- 167
x"01d00",-- 464
x"fb2e0",-- -1234
x"04fe0",-- 1278
x"fdd60",-- -554
x"00280",-- 40
x"07580",-- 1880
x"f9df0",-- -1569
x"fd440",-- -700
x"05220",-- 1314
x"007a0",-- 122
x"ffdf0",-- -33
x"fe8f0",-- -369
x"fa080",-- -1528
x"03d10",-- 977
x"01f10",-- 497
x"fec10",-- -319
x"014f0",-- 335
x"fcb90",-- -839
x"00280",-- 40
x"06860",-- 1670
x"fc0d0",-- -1011
x"fd3f0",-- -705
x"04550",-- 1109
x"fc370",-- -969
x"fd2e0",-- -722
x"04ac0",-- 1196
x"feda0",-- -294
x"00320",-- 50
x"01440",-- 324
x"f9f40",-- -1548
x"03900",-- 912
x"06890",-- 1673
x"fa3e0",-- -1474
x"fe960",-- -362
x"03d50",-- 981
x"01120",-- 274
x"04490",-- 1097
x"fe7b0",-- -389
x"faf00",-- -1296
x"053a0",-- 1338
x"01e20",-- 482
x"ff470",-- -185
x"03040",-- 772
x"fdfd0",-- -515
x"fbbd0",-- -1091
x"00690",-- 105
x"02690",-- 617
x"01ae0",-- 430
x"fca30",-- -861
x"fbe50",-- -1051
x"03e70",-- 999
x"01470",-- 327
x"fdab0",-- -597
x"fee30",-- -285
x"fea80",-- -344
x"025a0",-- 602
x"fe710",-- -399
x"fc6e0",-- -914
x"03fe0",-- 1022
x"00ad0",-- 173
x"fd2e0",-- -722
x"03290",-- 809
x"04530",-- 1107
x"fd9c0",-- -612
x"fe8a0",-- -374
x"01e50",-- 485
x"03df0",-- 991
x"ffea0",-- -22
x"ff600",-- -160
x"007a0",-- 122
x"fd110",-- -751
x"00410",-- 65
x"ff6a0",-- -150
x"fe280",-- -472
x"045c0",-- 1116
x"01d00",-- 464
x"fd040",-- -764
x"00780",-- 120
x"00b90",-- 185
x"fd830",-- -637
x"019a0",-- 410
x"01bd0",-- 445
x"fd330",-- -717
x"01030",-- 259
x"fbe00",-- -1056
x"ff3d0",-- -195
x"06730",-- 1651
x"f8260",-- -2010
x"ff580",-- -168
x"05120",-- 1298
x"fd330",-- -717
x"fea50",-- -347
x"03a60",-- 934
x"00490",-- 73
x"fdcb0",-- -565
x"01470",-- 327
x"fd3a0",-- -710
x"04700",-- 1136
x"01440",-- 324
x"fa6b0",-- -1429
x"05f30",-- 1523
x"014f0",-- 335
x"fa050",-- -1531
x"00e90",-- 233
x"01d80",-- 472
x"fdea0",-- -534
x"00350",-- 53
x"00250",-- 37
x"fe890",-- -375
x"ffd10",-- -47
x"fcd20",-- -814
x"ff670",-- -153
x"03e20",-- 994
x"fe760",-- -394
x"fe5a0",-- -422
x"02500",-- 592
x"fedf0",-- -289
x"fd070",-- -761
x"03040",-- 772
x"02990",-- 665
x"fe890",-- -375
x"fe5a0",-- -422
x"fe850",-- -379
x"03a90",-- 937
x"ffc90",-- -55
x"fd860",-- -634
x"010d0",-- 269
x"02030",-- 515
x"fc5c0",-- -932
x"006e0",-- 110
x"02ca0",-- 714
x"fe9b0",-- -357
x"fe0c0",-- -500
x"00520",-- 82
x"03790",-- 889
x"ffcc0",-- -52
x"fe0d0",-- -499
x"00230",-- 35
x"022b0",-- 555
x"003a0",-- 58
x"01240",-- 292
x"01560",-- 342
x"ff710",-- -143
x"fe730",-- -397
x"ff9e0",-- -98
x"017b0",-- 379
x"01ba0",-- 442
x"fe490",-- -439
x"fedc0",-- -292
x"03450",-- 837
x"00620",-- 98
x"fe070",-- -505
x"01e90",-- 489
x"feac0",-- -340
x"fd470",-- -697
x"02410",-- 577
x"fd040",-- -764
x"fd4c0",-- -692
x"00d00",-- 208
x"ff6a0",-- -150
x"020f0",-- 527
x"fff30",-- -13
x"ff860",-- -122
x"fd2f0",-- -721
x"ff8b0",-- -117
x"02640",-- 612
x"00700",-- 112
x"fffb0",-- -5
x"002b0",-- 43
x"ff300",-- -208
x"ffb50",-- -75
x"032b0",-- 811
x"00cb0",-- 203
x"fe2b0",-- -469
x"01580",-- 344
x"00fc0",-- 252
x"00f50",-- 245
x"02200",-- 544
x"ff3a0",-- -198
x"fff40",-- -12
x"00070",-- 7
x"ff900",-- -112
x"fffd0",-- -3
x"fc9e0",-- -866
x"fcf00",-- -784
x"fd270",-- -729
x"00960",-- 150
x"023f0",-- 575
x"fc230",-- -989
x"fdb50",-- -587
x"00a70",-- 167
x"ffd60",-- -42
x"00a30",-- 163
x"00190",-- 25
x"fee40",-- -284
x"ff2c0",-- -212
x"031d0",-- 797
x"01440",-- 324
x"fda40",-- -604
x"ff920",-- -110
x"02640",-- 612
x"01970",-- 407
x"ff7c0",-- -132
x"012c0",-- 300
x"00610",-- 97
x"fec50",-- -315
x"fec50",-- -315
x"01290",-- 297
x"ff5d0",-- -163
x"fe3f0",-- -449
x"01bc0",-- 444
x"023c0",-- 572
x"ffbc0",-- -68
x"fd830",-- -637
x"fd510",-- -687
x"00a30",-- 163
x"00980",-- 152
x"fe610",-- -415
x"030d0",-- 781
x"ff850",-- -123
x"fcad0",-- -851
x"01400",-- 320
x"01580",-- 344
x"00fe0",-- 254
x"03450",-- 837
x"00430",-- 67
x"fed90",-- -295
x"00ff0",-- 255
x"01970",-- 407
x"02210",-- 545
x"ff240",-- -220
x"ff2e0",-- -210
x"00960",-- 150
x"00ef0",-- 239
x"ffa30",-- -93
x"008f0",-- 143
x"ffab0",-- -85
x"fcc60",-- -826
x"00320",-- 50
x"01810",-- 385
x"ff040",-- -252
x"00230",-- 35
x"ffdf0",-- -33
x"fefd0",-- -259
x"00a70",-- 167
x"01150",-- 277
x"ffd10",-- -47
x"ff1f0",-- -225
x"ff270",-- -217
x"fe800",-- -384
x"01a10",-- 417
x"018a0",-- 394
x"feac0",-- -340
x"00f00",-- 240
x"01ad0",-- 429
x"ff290",-- -215
x"ff6f0",-- -145
x"012e0",-- 302
x"00490",-- 73
x"ff3d0",-- -195
x"ff5d0",-- -163
x"01c20",-- 450
x"004e0",-- 78
x"fdf10",-- -527
x"00d50",-- 213
x"fee30",-- -285
x"ffd50",-- -43
x"02a30",-- 675
x"00ed0",-- 237
x"00120",-- 18
x"01510",-- 337
x"01d30",-- 467
x"fe610",-- -415
x"fee80",-- -280
x"01fd0",-- 509
x"00fa0",-- 250
x"ff0e0",-- -242
x"fd5b0",-- -677
x"fe730",-- -397
x"fff40",-- -12
x"016d0",-- 365
x"00cf0",-- 207
x"fc980",-- -872
x"fccd0",-- -819
x"00fc0",-- 252
x"01fe0",-- 510
x"003a0",-- 58
x"ff220",-- -222
x"fe690",-- -407
x"00570",-- 87
x"04620",-- 1122
x"03bd0",-- 957
x"fe3e0",-- -450
x"fcd70",-- -809
x"fede0",-- -290
x"02fe0",-- 766
x"04660",-- 1126
x"00000",-- 0
x"fd5d0",-- -675
x"fdf90",-- -519
x"00210",-- 33
x"01100",-- 272
x"ffba0",-- -70
x"fce60",-- -794
x"fc5f0",-- -929
x"fe620",-- -414
x"00ed0",-- 237
x"012e0",-- 302
x"fdf60",-- -522
x"fb620",-- -1182
x"fcca0",-- -822
x"fe690",-- -407
x"00fe0",-- 254
x"02c30",-- 707
x"ff620",-- -158
x"fe8f0",-- -369
x"ff350",-- -203
x"00030",-- 3
x"fefd0",-- -259
x"000d0",-- 13
x"021c0",-- 540
x"ff580",-- -168
x"ff2e0",-- -210
x"00730",-- 115
x"00840",-- 132
x"ff990",-- -103
x"ff4c0",-- -180
x"02690",-- 617
x"00cf0",-- 207
x"fa430",-- -1469
x"fd2e0",-- -722
x"01100",-- 272
x"00bb0",-- 187
x"00690",-- 105
x"fe4d0",-- -435
x"ffcc0",-- -52
x"004d0",-- 77
x"01740",-- 372
x"02430",-- 579
x"01450",-- 325
x"00b90",-- 185
x"fe8f0",-- -369
x"ffda0",-- -38
x"03260",-- 806
x"02ad0",-- 685
x"ff630",-- -157
x"00640",-- 100
x"026e0",-- 622
x"003a0",-- 58
x"fee10",-- -287
x"00f50",-- 245
x"00280",-- 40
x"fe7d0",-- -387
x"ffc10",-- -63
x"009b0",-- 155
x"021b0",-- 539
x"000d0",-- 13
x"fdec0",-- -532
x"fe6b0",-- -405
x"fe0a0",-- -502
x"ffba0",-- -70
x"02d10",-- 721
x"02160",-- 534
x"ff270",-- -217
x"00020",-- 2
x"02f20",-- 754
x"02430",-- 579
x"ffbd0",-- -67
x"000a0",-- 10
x"00530",-- 83
x"01bf0",-- 447
x"02170",-- 535
x"00670",-- 103
x"ff2b0",-- -213
x"fee60",-- -282
x"fe9e0",-- -354
x"ffb20",-- -78
x"01060",-- 262
x"fefc0",-- -260
x"fd670",-- -665
x"ff420",-- -190
x"00580",-- 88
x"ffd50",-- -43
x"fe500",-- -432
x"fdbd0",-- -579
x"fee60",-- -282
x"ffa90",-- -87
x"02580",-- 600
x"03650",-- 869
x"01540",-- 340
x"ffd60",-- -42
x"fec60",-- -314
x"00050",-- 5
x"00210",-- 33
x"003a0",-- 58
x"01fd0",-- 509
x"01ad0",-- 429
x"ffa30",-- -93
x"ff830",-- -125
x"00e60",-- 230
x"00ef0",-- 239
x"00e10",-- 225
x"00730",-- 115
x"ff1d0",-- -227
x"ffb20",-- -78
x"00cf0",-- 207
x"01180",-- 280
x"00700",-- 112
x"ffd50",-- -43
x"00190",-- 25
x"00f40",-- 244
x"00440",-- 68
x"feda0",-- -294
x"fec10",-- -319
x"fea00",-- -352
x"ffa40",-- -92
x"01880",-- 392
x"02910",-- 657
x"ff110",-- -239
x"fc620",-- -926
x"ff100",-- -240
x"00760",-- 118
x"01b50",-- 437
x"01150",-- 277
x"fdf30",-- -525
x"fd8b0",-- -629
x"ffce0",-- -50
x"ff970",-- -105
x"ff1f0",-- -225
x"000c0",-- 12
x"fe370",-- -457
x"fe850",-- -379
x"024b0",-- 587
x"01710",-- 369
x"fd990",-- -615
x"fd990",-- -615
x"ffb50",-- -75
x"00350",-- 53
x"002f0",-- 47
x"ff380",-- -200
x"fe7b0",-- -389
x"ffc20",-- -62
x"004e0",-- 78
x"01590",-- 345
x"00d50",-- 213
x"fd100",-- -752
x"fdfb0",-- -517
x"010d0",-- 269
x"00ed0",-- 237
x"fff10",-- -15
x"006b0",-- 107
x"ff2e0",-- -210
x"fd450",-- -699
x"fdbd0",-- -579
x"ff630",-- -157
x"01d50",-- 469
x"02500",-- 592
x"001c0",-- 28
x"fe6b0",-- -405
x"febb0",-- -325
x"ff800",-- -128
x"023a0",-- 570
x"03ab0",-- 939
x"00a00",-- 160
x"fe2a0",-- -470
x"fe660",-- -410
x"ffbc0",-- -68
x"02340",-- 564
x"039e0",-- 926
x"01490",-- 329
x"fdc40",-- -572
x"fdd30",-- -557
x"006b0",-- 107
x"01310",-- 305
x"01090",-- 265
x"00c00",-- 192
x"00cd0",-- 205
x"00b20",-- 178
x"00670",-- 103
x"006e0",-- 110
x"002d0",-- 45
x"00a30",-- 163
x"00430",-- 67
x"01620",-- 354
x"02bc0",-- 700
x"000d0",-- 13
x"fe340",-- -460
x"001b0",-- 27
x"02cc0",-- 716
x"03490",-- 841
x"00e90",-- 233
x"00160",-- 22
x"02120",-- 530
x"037b0",-- 891
x"03950",-- 917
x"03100",-- 784
x"00b10",-- 177
x"fefd0",-- -259
x"00730",-- 115
x"02d90",-- 729
x"046c0",-- 1132
x"04480",-- 1096
x"010b0",-- 267
x"fd1f0",-- -737
x"ff860",-- -122
x"01f90",-- 505
x"023e0",-- 574
x"02ca0",-- 714
x"01180",-- 280
x"00020",-- 2
x"00430",-- 67
x"ffa60",-- -90
x"ff800",-- -128
x"012e0",-- 302
x"01ee0",-- 494
x"ffbf0",-- -65
x"ffb70",-- -73
x"ffa60",-- -90
x"00170",-- 23
x"02320",-- 562
x"00c10",-- 193
x"fdad0",-- -595
x"fdd10",-- -559
x"ffa40",-- -92
x"01510",-- 337
x"01bf0",-- 447
x"feb20",-- -334
x"fbe00",-- -1056
x"fbe00",-- -1056
x"fbad0",-- -1107
x"fccd0",-- -819
x"ff110",-- -239
x"fdc40",-- -572
x"fb970",-- -1129
x"fb6c0",-- -1172
x"fb0b0",-- -1269
x"fab60",-- -1354
x"fae30",-- -1309
x"fab60",-- -1354
x"fac30",-- -1341
x"fc190",-- -999
x"fbae0",-- -1106
x"fac00",-- -1344
x"fb400",-- -1216
x"fc580",-- -936
x"fb360",-- -1226
x"fa980",-- -1384
x"fc340",-- -972
x"fcad0",-- -851
x"fbfd0",-- -1027
x"fae60",-- -1306
x"faa20",-- -1374
x"fc690",-- -919
x"fda80",-- -600
x"fdd00",-- -560
x"fd4f0",-- -689
x"fcd40",-- -812
x"fc550",-- -939
x"fc850",-- -891
x"fecd0",-- -307
x"ff1f0",-- -225
x"ff2b0",-- -213
x"00570",-- 87
x"000c0",-- 12
x"fede0",-- -290
x"fee90",-- -279
x"fec00",-- -320
x"fe070",-- -505
x"ffbd0",-- -67
x"01bc0",-- 444
x"03530",-- 851
x"032e0",-- 814
x"02a00",-- 672
x"03da0",-- 986
x"03bd0",-- 957
x"02870",-- 647
x"039e0",-- 926
x"05600",-- 1376
x"05a40",-- 1444
x"056c0",-- 1388
x"04ef0",-- 1263
x"04230",-- 1059
x"04530",-- 1107
x"05400",-- 1344
x"06810",-- 1665
x"071f0",-- 1823
x"06620",-- 1634
x"05c40",-- 1476
x"06e60",-- 1766
x"082d0",-- 2093
x"09650",-- 2405
x"09e40",-- 2532
x"07900",-- 1936
x"05fb0",-- 1531
x"086b0",-- 2155
x"0bfb0",-- 3067
x"0c2f0",-- 3119
x"0acf0",-- 2767
x"0a680",-- 2664
x"09710",-- 2417
x"07c20",-- 1986
x"08c20",-- 2242
x"09330",-- 2355
x"07a40",-- 1956
x"06dc0",-- 1756
x"08910",-- 2193
x"09ec0",-- 2540
x"08e30",-- 2275
x"08340",-- 2100
x"08c50",-- 2245
x"082f0",-- 2095
x"03680",-- 872
x"feb20",-- -334
x"ffb70",-- -73
x"01900",-- 400
x"fedc0",-- -292
x"fa520",-- -1454
x"f90b0",-- -1781
x"f6e30",-- -2333
x"f35c0",-- -3236
x"eff20",-- -4110
x"ef9a0",-- -4198
x"f1020",-- -3838
x"f1240",-- -3804
x"f0cb0",-- -3893
x"eff20",-- -4110
x"ef290",-- -4311
x"f0cb0",-- -3893
x"f1d80",-- -3624
x"ef220",-- -4318
x"ed480",-- -4792
x"ef4a0",-- -4278
x"f3bd0",-- -3139
x"f6d00",-- -2352
x"f5200",-- -2784
x"f2cf0",-- -3377
x"f29b0",-- -3429
x"f4000",-- -3072
x"f7630",-- -2205
x"fa170",-- -1513
x"f95e0",-- -1698
x"f6760",-- -2442
x"f4cd0",-- -2867
x"f59d0",-- -2659
x"f7ad0",-- -2131
x"f8390",-- -1991
x"f61e0",-- -2530
x"f5950",-- -2667
x"f7fe0",-- -2050
x"f8e10",-- -1823
x"f9a60",-- -1626
x"f9d50",-- -1579
x"f8ff0",-- -1793
x"fa140",-- -1516
x"fd3d0",-- -707
x"feaf0",-- -337
x"fe8f0",-- -369
x"ffa30",-- -93
x"00f50",-- 245
x"02e10",-- 737
x"045f0",-- 1119
x"03fe0",-- 1022
x"04080",-- 1032
x"05c40",-- 1476
x"07e70",-- 2023
x"09d50",-- 2517
x"09a10",-- 2465
x"08b10",-- 2225
x"09920",-- 2450
x"0c2a0",-- 3114
x"0e410",-- 3649
x"0d600",-- 3424
x"0bb00",-- 2992
x"0b010",-- 2817
x"0b710",-- 2929
x"0c140",-- 3092
x"0dab0",-- 3499
x"0ea70",-- 3751
x"0d150",-- 3349
x"0d4e0",-- 3406
x"10640",-- 4196
x"12140",-- 4628
x"12200",-- 4640
x"10400",-- 4160
x"0f1f0",-- 3871
x"114a0",-- 4426
x"12190",-- 4633
x"12b90",-- 4793
x"137e0",-- 4990
x"13a10",-- 5025
x"10140",-- 4116
x"0e050",-- 3589
x"108b0",-- 4235
x"10fe0",-- 4350
x"0e280",-- 3624
x"0f8a0",-- 3978
x"106b0",-- 4203
x"0c910",-- 3217
x"063f0",-- 1599
x"04ed0",-- 1261
x"05e20",-- 1506
x"ff860",-- -122
x"faa30",-- -1373
x"f6cb0",-- -2357
x"f4870",-- -2937
x"f41c0",-- -3044
x"f2da0",-- -3366
x"f17e0",-- -3714
x"ee930",-- -4461
x"eb3d0",-- -5315
x"e95e0",-- -5794
x"ea460",-- -5562
x"eb430",-- -5309
x"e86a0",-- -6038
x"e5cf0",-- -6705
x"e46c0",-- -7060
x"e7830",-- -6269
x"ef700",-- -4240
x"f1fe0",-- -3586
x"efea0",-- -4118
x"ece90",-- -4887
x"eda20",-- -4702
x"f1ca0",-- -3638
x"f64e0",-- -2482
x"f7470",-- -2233
x"f4bb0",-- -2885
x"f3dd0",-- -3107
x"f3c50",-- -3131
x"f44d0",-- -2995
x"f51f0",-- -2785
x"f4500",-- -2992
x"f2c00",-- -3392
x"f2640",-- -3484
x"f2ac0",-- -3412
x"f4700",-- -2960
x"f4940",-- -2924
x"f3f30",-- -3085
x"f4070",-- -3065
x"f4a80",-- -2904
x"f6eb0",-- -2325
x"f9570",-- -1705
x"fa210",-- -1503
x"fa7a0",-- -1414
x"fc430",-- -957
x"fe730",-- -397
x"ffd00",-- -48
x"00b90",-- 185
x"01990",-- 409
x"04a50",-- 1189
x"08440",-- 2116
x"09530",-- 2387
x"09d50",-- 2517
x"0a320",-- 2610
x"09e00",-- 2528
x"0ab60",-- 2742
x"0bcc0",-- 3020
x"0d3d0",-- 3389
x"0ed10",-- 3793
x"0ee00",-- 3808
x"0e4b0",-- 3659
x"0e340",-- 3636
x"0ef40",-- 3828
x"10ca0",-- 4298
x"13aa0",-- 5034
x"145c0",-- 5212
x"12e50",-- 4837
x"12570",-- 4695
x"13df0",-- 5087
x"16400",-- 5696
x"18890",-- 6281
x"19560",-- 6486
x"19710",-- 6513
x"18730",-- 6259
x"17e70",-- 6119
x"19080",-- 6408
x"17120",-- 5906
x"160c0",-- 5644
x"186d0",-- 6253
x"1ba30",-- 7075
x"1e220",-- 7714
x"1c8e0",-- 7310
x"1a4f0",-- 6735
x"15d70",-- 5591
x"0f950",-- 3989
x"06190",-- 1561
x"00120",-- 18
x"fec60",-- -314
x"fb3e0",-- -1218
x"f7020",-- -2302
x"f5d30",-- -2605
x"f06b0",-- -3989
x"e8790",-- -6023
x"e6d80",-- -6440
x"e9420",-- -5822
x"e8850",-- -6011
x"e5cc0",-- -6708
x"e80b0",-- -6133
x"ea510",-- -5551
x"eb1b0",-- -5349
x"ec240",-- -5084
x"ebd60",-- -5162
x"eafc0",-- -5380
x"ee210",-- -4575
x"f1ae0",-- -3666
x"f1930",-- -3693
x"f1de0",-- -3618
x"f3ef0",-- -3089
x"f26b0",-- -3477
x"f04b0",-- -4021
x"f1b60",-- -3658
x"f0700",-- -3984
x"ef160",-- -4330
x"f0710",-- -3983
x"f06e0",-- -3986
x"ee2e0",-- -4562
x"ebbb0",-- -5189
x"eade0",-- -5410
x"eabe0",-- -5442
x"ec2d0",-- -5075
x"ef5c0",-- -4260
x"efdd0",-- -4131
x"f0320",-- -4046
x"f1590",-- -3751
x"f2b60",-- -3402
x"f4ad0",-- -2899
x"f6710",-- -2447
x"f8e30",-- -1821
x"f9720",-- -1678
x"fb2c0",-- -1236
x"fc980",-- -872
x"fca80",-- -856
x"fe250",-- -475
x"00c30",-- 195
x"02200",-- 544
x"03d60",-- 982
x"04f00",-- 1264
x"04fa0",-- 1274
x"058f0",-- 1423
x"07940",-- 1940
x"09030",-- 2307
x"0a7a0",-- 2682
x"0c1b0",-- 3099
x"0cb80",-- 3256
x"0cff0",-- 3327
x"0d790",-- 3449
x"0f630",-- 3939
x"10fa0",-- 4346
x"10ef0",-- 4335
x"11e60",-- 4582
x"14890",-- 5257
x"15240",-- 5412
x"157e0",-- 5502
x"162c0",-- 5676
x"18730",-- 6259
x"19f80",-- 6648
x"1bfa0",-- 7162
x"1db90",-- 7609
x"1c680",-- 7272
x"1d4e0",-- 7502
x"215a0",-- 8538
x"26700",-- 9840
x"24d90",-- 9433
x"1b1a0",-- 6938
x"19e90",-- 6633
x"21f00",-- 8688
x"2a2f0",-- 10799
x"25cb0",-- 9675
x"11130",-- 4371
x"ffe90",-- -23
x"f8a30",-- -1885
x"fe6b0",-- -405
x"ff110",-- -239
x"f6aa0",-- -2390
x"ee280",-- -4568
x"e5cf0",-- -6705
x"e2910",-- -7535
x"e3ba0",-- -7238
x"e71b0",-- -6373
x"e44b0",-- -7093
x"dd160",-- -8938
x"df4d0",-- -8371
x"e9830",-- -5757
x"ef090",-- -4343
x"f2170",-- -3561
x"f02d0",-- -4051
x"f1020",-- -3838
x"f4e90",-- -2839
x"fac10",-- -1343
x"fe6c0",-- -404
x"fbf60",-- -1034
x"fb5c0",-- -1188
x"fa660",-- -1434
x"fabc0",-- -1348
x"f97c0",-- -1668
x"f5b60",-- -2634
x"f1200",-- -3808
x"ed3e0",-- -4802
x"eb560",-- -5290
x"ea780",-- -5512
x"e5cf0",-- -6705
x"e3000",-- -7424
x"e31d0",-- -7395
x"e7cf0",-- -6193
x"ebd40",-- -5164
x"ec850",-- -4987
x"ee190",-- -4583
x"ed7f0",-- -4737
x"f0030",-- -4093
x"f4b20",-- -2894
x"f9e90",-- -1559
x"fc610",-- -927
x"fc9e0",-- -866
x"fe2d0",-- -467
x"ffea0",-- -22
x"00a20",-- 162
x"01e90",-- 489
x"01580",-- 344
x"018b0",-- 395
x"02f70",-- 759
x"04300",-- 1072
x"051d0",-- 1309
x"03e00",-- 992
x"036f0",-- 879
x"034c0",-- 844
x"05530",-- 1363
x"07720",-- 1906
x"08580",-- 2136
x"08340",-- 2100
x"08dc0",-- 2268
x"0b600",-- 2912
x"0eae0",-- 3758
x"10cd0",-- 4301
x"12f00",-- 4848
x"14cf0",-- 5327
x"16280",-- 5672
x"183c0",-- 6204
x"19030",-- 6403
x"1a410",-- 6721
x"1acd0",-- 6861
x"1c590",-- 7257
x"1cb80",-- 7352
x"1e180",-- 7704
x"20b00",-- 8368
x"25100",-- 9488
x"287a0",-- 10362
x"2a240",-- 10788
x"27e80",-- 10216
x"25c10",-- 9665
x"25ce0",-- 9678
x"24b60",-- 9398
x"1a6e0",-- 6766
x"07c90",-- 1993
x"f9660",-- -1690
x"f6990",-- -2407
x"fa430",-- -1469
x"f7970",-- -2153
x"eee80",-- -4376
x"e19a0",-- -7782
x"db720",-- -9358
x"da0f0",-- -9713
x"dda70",-- -8793
x"df360",-- -8394
x"dd370",-- -8905
x"e02b0",-- -8149
x"e5e20",-- -6686
x"ef9c0",-- -4196
x"f6b40",-- -2380
x"f8b90",-- -1863
x"f8ff0",-- -1793
x"fb480",-- -1208
x"014a0",-- 330
x"07fd0",-- 2045
x"09560",-- 2390
x"08db0",-- 2267
x"04ae0",-- 1198
x"015d0",-- 349
x"fdd60",-- -554
x"f9880",-- -1656
x"f5060",-- -2810
x"ee8a0",-- -4470
x"eaa80",-- -5464
x"e7470",-- -6329
x"e42d0",-- -7123
x"e0f00",-- -7952
x"dfac0",-- -8276
x"e1a90",-- -7767
x"e5fb0",-- -6661
x"ea6e0",-- -5522
x"edc40",-- -4668
x"ef5b0",-- -4261
x"f2280",-- -3544
x"f56f0",-- -2705
x"f86e0",-- -1938
x"f9560",-- -1706
x"fb240",-- -1244
x"ff540",-- -172
x"038f0",-- 911
x"04850",-- 1157
x"022b0",-- 555
x"001e0",-- 30
x"ff6d0",-- -147
x"01600",-- 352
x"03440",-- 836
x"033d0",-- 829
x"00aa0",-- 170
x"fe730",-- -397
x"feca0",-- -310
x"00b70",-- 183
x"02730",-- 627
x"02e00",-- 736
x"02710",-- 625
x"033f0",-- 831
x"05dd0",-- 1501
x"088c0",-- 2188
x"0b2b0",-- 2859
x"0c750",-- 3189
x"0eed0",-- 3821
x"11a10",-- 4513
x"16480",-- 5704
x"187f0",-- 6271
x"19330",-- 6451
x"19ab0",-- 6571
x"1b5b0",-- 7003
x"1c980",-- 7320
x"1c400",-- 7232
x"1ddc0",-- 7644
x"1dd50",-- 7637
x"21710",-- 8561
x"24c70",-- 9415
x"29ba0",-- 10682
x"29b00",-- 10672
x"28fb0",-- 10491
x"2c700",-- 11376
x"2d350",-- 11573
x"23da0",-- 9178
x"0cf00",-- 3312
x"f2930",-- -3437
x"e92a0",-- -5846
x"ece60",-- -4890
x"f3040",-- -3324
x"f1560",-- -3754
x"e7ca0",-- -6198
x"de4e0",-- -8626
x"d22c0",-- -11732
x"d2170",-- -11753
x"d8790",-- -10119
x"dd0a0",-- -8950
x"df360",-- -8394
x"e4530",-- -7085
x"ef900",-- -4208
x"f7ae0",-- -2130
x"fb9a0",-- -1126
x"fdce0",-- -562
x"ff060",-- -250
x"03880",-- 904
x"0bf10",-- 3057
x"12e30",-- 4835
x"142c0",-- 5164
x"0c930",-- 3219
x"06de0",-- 1758
x"031f0",-- 799
x"01620",-- 354
x"fb3e0",-- -1218
x"f2760",-- -3466
x"ebfc0",-- -5124
x"e69b0",-- -6501
x"e2b70",-- -7497
x"df130",-- -8429
x"dcf80",-- -8968
x"dde30",-- -8733
x"e0c80",-- -7992
x"e6c10",-- -6463
x"ec470",-- -5049
x"efd80",-- -4136
x"ef570",-- -4265
x"eec10",-- -4415
x"f6f50",-- -2315
x"01260",-- 294
x"07d30",-- 2003
x"06a90",-- 1705
x"03ba0",-- 954
x"003e0",-- 62
x"fdbd0",-- -579
x"00960",-- 150
x"02a80",-- 680
x"03490",-- 841
x"022a0",-- 554
x"00ef0",-- 239
x"ff400",-- -192
x"fce90",-- -791
x"fb8a0",-- -1142
x"fa460",-- -1466
x"fa670",-- -1433
x"fd440",-- -700
x"ff9a0",-- -102
x"01260",-- 294
x"00da0",-- 218
x"018f0",-- 399
x"03900",-- 912
x"063e0",-- 1598
x"0a140",-- 2580
x"0c5a0",-- 3162
x"0fb00",-- 4016
x"11a60",-- 4518
x"12f50",-- 4853
x"13770",-- 4983
x"147a0",-- 5242
x"17460",-- 5958
x"1a950",-- 6805
x"1c7f0",-- 7295
x"1b3d0",-- 6973
x"18340",-- 6196
x"178f0",-- 6031
x"1a840",-- 6788
x"1fdf0",-- 8159
x"24510",-- 9297
x"25a00",-- 9632
x"27830",-- 10115
x"29e80",-- 10728
x"2e570",-- 11863
x"2bfc0",-- 11260
x"1c550",-- 7253
x"fe230",-- -477
x"e6370",-- -6601
x"e4a10",-- -7007
x"edb80",-- -4680
x"f1bf0",-- -3649
x"ec050",-- -5115
x"e5de0",-- -6690
x"df140",-- -8428
x"d9220",-- -9950
x"da030",-- -9725
x"ddce0",-- -8754
x"e3250",-- -7387
x"eb4d0",-- -5299
x"f5bd0",-- -2627
x"00bc0",-- 188
x"052e0",-- 1326
x"05040",-- 1284
x"03310",-- 817
x"04430",-- 1091
x"0b560",-- 2902
x"113d0",-- 4413
x"10f90",-- 4345
x"0a900",-- 2704
x"050b0",-- 1291
x"01810",-- 385
x"f9a10",-- -1631
x"edca0",-- -4662
x"e5a60",-- -6746
x"e3250",-- -7387
x"e2260",-- -7642
x"ddca0",-- -8758
x"dbc70",-- -9273
x"dbd60",-- -9258
x"dcda0",-- -8998
x"e2c80",-- -7480
x"eb790",-- -5255
x"f3d60",-- -3114
x"f7fe0",-- -2050
x"fb420",-- -1214
x"fefa0",-- -262
x"01a10",-- 417
x"04ac0",-- 1196
x"06190",-- 1561
x"05fe0",-- 1534
x"03c70",-- 967
x"02050",-- 517
x"02580",-- 600
x"01670",-- 359
x"ff150",-- -235
x"fa160",-- -1514
x"f8a20",-- -1886
x"f7970",-- -2153
x"f4850",-- -2939
x"f3a90",-- -3159
x"f3a70",-- -3161
x"f75b0",-- -2213
x"fa1b0",-- -1509
x"fcd70",-- -809
x"fff60",-- -10
x"01da0",-- 474
x"05990",-- 1433
x"085c0",-- 2140
x"0b010",-- 2817
x"0d580",-- 3416
x"0d270",-- 3367
x"0da60",-- 3494
x"0dd30",-- 3539
x"0e900",-- 3728
x"0d9c0",-- 3484
x"0b1c0",-- 2844
x"0a430",-- 2627
x"09900",-- 2448
x"0bae0",-- 2990
x"0cb30",-- 3251
x"0cf00",-- 3312
x"0e370",-- 3639
x"11530",-- 4435
x"154f0",-- 5455
x"17f10",-- 6129
x"19c60",-- 6598
x"1cea0",-- 7402
x"21d70",-- 8663
x"28cf0",-- 10447
x"2fde0",-- 12254
x"335d0",-- 13149
x"32c50",-- 12997
x"2fcb0",-- 12235
x"28de0",-- 10462
x"13dc0",-- 5084
x"f65f0",-- -2465
x"e2f60",-- -7434
x"e3c70",-- -7225
x"ec820",-- -4990
x"ec7e0",-- -4994
x"e57c0",-- -6788
x"dd840",-- -8828
x"d5130",-- -10989
x"d27b0",-- -11653
x"d6650",-- -10651
x"dfd10",-- -8239
x"e95b0",-- -5797
x"f13e0",-- -3778
x"fddf0",-- -545
x"07f90",-- 2041
x"0d150",-- 3349
x"0c340",-- 3124
x"0ae80",-- 2792
x"0e4d0",-- 3661
x"13ff0",-- 5119
x"18de0",-- 6366
x"180e0",-- 6158
x"10cc0",-- 4300
x"05800",-- 1408
x"f92f0",-- -1745
x"f0480",-- -4024
x"e8d20",-- -5934
x"de6a0",-- -8598
x"d5c80",-- -10808
x"d3c20",-- -11326
x"d7950",-- -10347
x"d8230",-- -10205
x"d7a90",-- -10327
x"daba0",-- -9542
x"e12c0",-- -7892
x"ea940",-- -5484
x"f4d50",-- -2859
x"fd9a0",-- -614
x"016f0",-- 367
x"03b30",-- 947
x"08700",-- 2160
x"0c340",-- 3124
x"0e5e0",-- 3678
x"0d6c0",-- 3436
x"0a120",-- 2578
x"04f40",-- 1268
x"ff5b0",-- -165
x"ff0b0",-- -245
x"fe2f0",-- -465
x"fd600",-- -672
x"f77a0",-- -2182
x"f0a50",-- -3931
x"ee800",-- -4480
x"ef5b0",-- -4261
x"f4530",-- -2989
x"f6940",-- -2412
x"f7340",-- -2252
x"f7db0",-- -2085
x"fbe00",-- -1056
x"03470",-- 839
x"08ca0",-- 2250
x"0b3d0",-- 2877
x"0bc90",-- 3017
x"0b0b0",-- 2827
x"0ca40",-- 3236
x"0e860",-- 3718
x"100a0",-- 4106
x"0f7e0",-- 3966
x"0df50",-- 3573
x"0dbf0",-- 3519
x"0c870",-- 3207
x"0d670",-- 3431
x"0d4e0",-- 3406
x"0dc10",-- 3521
x"0f8f0",-- 3983
x"14320",-- 5170
x"186b0",-- 6251
x"1a430",-- 6723
x"194c0",-- 6476
x"18890",-- 6281
x"1bc90",-- 7113
x"212b0",-- 8491
x"2a860",-- 10886
x"30430",-- 12355
x"33e60",-- 13286
x"337d0",-- 13181
x"29ad0",-- 10669
x"13360",-- 4918
x"f34c0",-- -3252
x"debe0",-- -8514
x"de470",-- -8633
x"e9a20",-- -5726
x"f04b0",-- -4021
x"ed970",-- -4713
x"e4c10",-- -6975
x"d9250",-- -9947
x"d34b0",-- -11445
x"d8a10",-- -10079
x"e2730",-- -7565
x"ebf90",-- -5127
x"f77f0",-- -2177
x"05ab0",-- 1451
x"0f5b0",-- 3931
x"0fd70",-- 4055
x"0d850",-- 3461
x"0a6b0",-- 2667
x"0ab60",-- 2742
x"0f9c0",-- 3996
x"15380",-- 5432
x"16410",-- 5697
x"0f220",-- 3874
x"056c0",-- 1388
x"f9ef0",-- -1553
x"ecd50",-- -4907
x"e1c20",-- -7742
x"dc210",-- -9183
x"dcbf0",-- -9025
x"d7be0",-- -10306
x"d12c0",-- -11988
x"d2420",-- -11710
x"d8ee0",-- -10002
x"e0530",-- -8109
x"e5900",-- -6768
x"eef00",-- -4368
x"f77a0",-- -2182
x"fdb50",-- -587
x"05ec0",-- 1516
x"0a910",-- 2705
x"0aaa0",-- 2730
x"0a050",-- 2565
x"0b970",-- 2967
x"0d0b0",-- 3339
x"0ae50",-- 2789
x"07630",-- 1891
x"00c30",-- 195
x"f8850",-- -1915
x"f2d20",-- -3374
x"f2e40",-- -3356
x"f40c0",-- -3060
x"f4e80",-- -2840
x"f4520",-- -2990
x"f0f00",-- -3856
x"f0660",-- -3994
x"f18e0",-- -3698
x"f6320",-- -2510
x"fb4f0",-- -1201
x"ffe90",-- -23
x"045f0",-- 1119
x"086e0",-- 2158
x"0bab0",-- 2987
x"0d300",-- 3376
x"0ca40",-- 3236
x"0c9a0",-- 3226
x"0d240",-- 3364
x"0e770",-- 3703
x"0f770",-- 3959
x"0e730",-- 3699
x"0cc70",-- 3271
x"0a370",-- 2615
x"09ae0",-- 2478
x"0ab60",-- 2742
x"0c5c0",-- 3164
x"0c7f0",-- 3199
x"0e250",-- 3621
x"12c00",-- 4800
x"16e60",-- 5862
x"1a140",-- 6676
x"1ac30",-- 6851
x"1a9a0",-- 6810
x"1d3a0",-- 7482
x"249c0",-- 9372
x"2f910",-- 12177
x"34bf0",-- 13503
x"36240",-- 13860
x"30f70",-- 12535
x"1dfb0",-- 7675
x"fdd10",-- -559
x"e1ef0",-- -7697
x"ddba0",-- -8774
x"e5790",-- -6791
x"ebfc0",-- -5124
x"eddb0",-- -4645
x"ea5f0",-- -5537
x"e0780",-- -8072
x"d64c0",-- -10676
x"d8740",-- -10124
x"e1f40",-- -7692
x"e9ea0",-- -5654
x"f55b0",-- -2725
x"03ec0",-- 1004
x"0f540",-- 3924
x"10e80",-- 4328
x"0f860",-- 3974
x"0de20",-- 3554
x"09ad0",-- 2477
x"0a700",-- 2672
x"0f710",-- 3953
x"13120",-- 4882
x"0f350",-- 3893
x"06a70",-- 1703
x"fc9b0",-- -869
x"efce0",-- -4146
x"e3180",-- -7400
x"db2c0",-- -9428
x"d91b0",-- -9957
x"dac80",-- -9528
x"da290",-- -9687
x"d7d10",-- -10287
x"d5ef0",-- -10769
x"db9b0",-- -9317
x"e7930",-- -6253
x"f2a30",-- -3421
x"fab20",-- -1358
x"fe9e0",-- -354
x"03540",-- 852
x"06960",-- 1686
x"09ea0",-- 2538
x"0af20",-- 2802
x"095e0",-- 2398
x"07940",-- 1940
x"063a0",-- 1594
x"04f20",-- 1266
x"00f50",-- 245
x"fadf0",-- -1313
x"f5400",-- -2752
x"f0760",-- -3978
x"ef420",-- -4286
x"f1a90",-- -3671
x"f4f30",-- -2829
x"f6b90",-- -2375
x"f4870",-- -2937
x"f4140",-- -3052
x"f47a0",-- -2950
x"f8cb0",-- -1845
x"fe7b0",-- -389
x"06250",-- 1573
x"0abe0",-- 2750
x"0edc0",-- 3804
x"11100",-- 4368
x"08580",-- 2136
x"09790",-- 2425
x"0d380",-- 3384
x"0ca40",-- 3236
x"0d2b0",-- 3371
x"09bc0",-- 2492
x"08db0",-- 2267
x"0a050",-- 2565
x"08c50",-- 2245
x"081b0",-- 2075
x"098a0",-- 2442
x"0a8e0",-- 2702
x"09f40",-- 2548
x"0e640",-- 3684
x"15300",-- 5424
x"18720",-- 6258
x"1aa90",-- 6825
x"1c320",-- 7218
x"1de10",-- 7649
x"22c90",-- 8905
x"29e40",-- 10724
x"310a0",-- 12554
x"333e0",-- 13118
x"35320",-- 13618
x"2e660",-- 11878
x"164f0",-- 5711
x"f3f30",-- -3085
x"db0a0",-- -9462
x"d7980",-- -10344
x"df190",-- -8423
x"eada0",-- -5414
x"ee320",-- -4558
x"e7090",-- -6391
x"e01f0",-- -8161
x"d8a80",-- -10072
x"dff10",-- -8207
x"e7fc0",-- -6148
x"ec990",-- -4967
x"fd5d0",-- -675
x"0d6c0",-- 3436
x"16250",-- 5669
x"134c0",-- 4940
x"15420",-- 5442
x"0de90",-- 3561
x"097e0",-- 2430
x"05ae0",-- 1454
x"09f10",-- 2545
x"10690",-- 4201
x"0c020",-- 3074
x"fed40",-- -300
x"f5070",-- -2809
x"eba60",-- -5210
x"d7480",-- -10424
x"d89e0",-- -10082
x"d58b0",-- -10869
x"dbb30",-- -9293
x"de240",-- -8668
x"dd1e0",-- -8930
x"dde50",-- -8731
x"df340",-- -8396
x"ed150",-- -4843
x"f9f90",-- -1543
x"023c0",-- 572
x"02a70",-- 679
x"06c50",-- 1733
x"0b2b0",-- 2859
x"0a6e0",-- 2670
x"07b30",-- 1971
x"055e0",-- 1374
x"034a0",-- 842
x"01440",-- 324
x"fe500",-- -432
x"fdcc0",-- -564
x"f8800",-- -1920
x"f1b60",-- -3658
x"ed6a0",-- -4758
x"eecd0",-- -4403
x"f3200",-- -3296
x"f3b00",-- -3152
x"f6bb0",-- -2373
x"f6a00",-- -2400
x"f8730",-- -1933
x"fb020",-- -1278
x"ff020",-- -254
x"02f90",-- 761
x"05f10",-- 1521
x"0c2d0",-- 3117
x"0f1f0",-- 3871
x"0f9a0",-- 3994
x"0c8c0",-- 3212
x"09850",-- 2437
x"08490",-- 2121
x"07a60",-- 1958
x"08c70",-- 2247
x"058b0",-- 1419
x"0cef0",-- 3311
x"09e00",-- 2528
x"03010",-- 769
x"052c0",-- 1324
x"05e90",-- 1513
x"0c910",-- 3217
x"0e570",-- 3671
x"0f150",-- 3861
x"17e40",-- 6116
x"1bc90",-- 7113
x"1c2c0",-- 7212
x"1e040",-- 7684
x"209d0",-- 8349
x"269d0",-- 9885
x"29780",-- 10616
x"2f850",-- 12165
x"339e0",-- 13214
x"33da0",-- 13274
x"28de0",-- 10462
x"08a50",-- 2213
x"e5020",-- -6910
x"d4380",-- -11208
x"d8bc0",-- -10052
x"e1b00",-- -7760
x"e6f50",-- -6411
x"eb520",-- -5294
x"eaa80",-- -5464
x"e30a0",-- -7414
x"e0a30",-- -8029
x"e4260",-- -7130
x"ec6c0",-- -5012
x"f1950",-- -3691
x"01b70",-- 439
x"170b0",-- 5899
x"1c8c0",-- 7308
x"1aae0",-- 6830
x"12fe0",-- 4862
x"0c0a0",-- 3082
x"05a90",-- 1449
x"01e40",-- 484
x"05790",-- 1401
x"06e60",-- 1766
x"01e90",-- 489
x"f8fd0",-- -1795
x"ef340",-- -4300
x"e45a0",-- -7078
x"d6b70",-- -10569
x"d28d0",-- -11635
x"d7340",-- -10444
x"de410",-- -8639
x"e15f0",-- -7841
x"e2740",-- -7564
x"e6990",-- -6503
x"ed9d0",-- -4707
x"f6cd0",-- -2355
x"fd490",-- -695
x"01060",-- 262
x"04f50",-- 1269
x"091f0",-- 2335
x"0ab80",-- 2744
x"09880",-- 2440
x"06500",-- 1616
x"00bb0",-- 187
x"fb7b0",-- -1157
x"fa3c0",-- -1476
x"fb520",-- -1198
x"f9d80",-- -1576
x"f4df0",-- -2849
x"ef9c0",-- -4196
x"eeed0",-- -4371
x"f1a40",-- -3676
x"f35e0",-- -3234
x"f5570",-- -2729
x"f7d60",-- -2090
x"fa440",-- -1468
x"fc890",-- -887
x"ff560",-- -170
x"01b20",-- 434
x"03fe0",-- 1022
x"08050",-- 2053
x"0c020",-- 3074
x"0e780",-- 3704
x"0fc40",-- 4036
x"0d760",-- 3446
x"09150",-- 2325
x"05fb0",-- 1531
x"05240",-- 1316
x"05ec0",-- 1516
x"063e0",-- 1598
x"06140",-- 1556
x"06030",-- 1539
x"057b0",-- 1403
x"068c0",-- 1676
x"0a6e0",-- 2670
x"0c4d0",-- 3149
x"0da30",-- 3491
x"11f10",-- 4593
x"18a40",-- 6308
x"1e4b0",-- 7755
x"20ea0",-- 8426
x"21f10",-- 8689
x"22590",-- 8793
x"23280",-- 9000
x"27e80",-- 10216
x"2ed30",-- 11987
x"31000",-- 12544
x"2f2d0",-- 12077
x"21640",-- 8548
x"03bf0",-- 959
x"e2490",-- -7607
x"d07b0",-- -12165
x"d5690",-- -10903
x"dd930",-- -8813
x"e3970",-- -7273
x"ea7b0",-- -5509
x"ef510",-- -4271
x"ed630",-- -4765
x"ead40",-- -5420
x"ee230",-- -4573
x"f2230",-- -3549
x"f85d0",-- -1955
x"05590",-- 1369
x"14e30",-- 5347
x"1dc80",-- 7624
x"1c320",-- 7218
x"132b0",-- 4907
x"08c70",-- 2247
x"feb70",-- -329
x"fa020",-- -1534
x"f92f0",-- -1745
x"fb1b0",-- -1253
x"faaa0",-- -1366
x"f7790",-- -2183
x"ef480",-- -4280
x"e1ce0",-- -7730
x"d6440",-- -10684
x"d3550",-- -11435
x"da3d0",-- -9667
x"e0650",-- -8091
x"e57e0",-- -6786
x"ead90",-- -5415
x"f2550",-- -3499
x"f93b0",-- -1733
x"fcbe0",-- -834
x"fed20",-- -302
x"007a0",-- 122
x"03490",-- 841
x"07ad0",-- 1965
x"0a630",-- 2659
x"09db0",-- 2523
x"033a0",-- 826
x"fb7e0",-- -1154
x"f61b0",-- -2533
x"f44d0",-- -2995
x"f5860",-- -2682
x"f41e0",-- -3042
x"f42f0",-- -3025
x"f37a0",-- -3206
x"f2f80",-- -3336
x"f4a00",-- -2912
x"f6be0",-- -2370
x"f6170",-- -2537
x"f75c0",-- -2212
x"fb800",-- -1152
x"00000",-- 0
x"04620",-- 1122
x"06760",-- 1654
x"09420",-- 2370
x"0aef0",-- 2799
x"0bd30",-- 3027
x"0c7d0",-- 3197
x"0c130",-- 3091
x"09740",-- 2420
x"06ea0",-- 1770
x"04d60",-- 1238
x"03b80",-- 952
x"023e0",-- 574
x"01740",-- 372
x"02640",-- 612
x"03e90",-- 1001
x"06c70",-- 1735
x"08930",-- 2195
x"0b650",-- 2917
x"0d1f0",-- 3359
x"0fba0",-- 4026
x"12dc0",-- 4828
x"17b20",-- 6066
x"1d9e0",-- 7582
x"20310",-- 8241
x"21b70",-- 8631
x"22540",-- 8788
x"24230",-- 9251
x"290d0",-- 10509
x"2db70",-- 11703
x"2dda0",-- 11738
x"2a8d0",-- 10893
x"1ef90",-- 7929
x"08bb0",-- 2235
x"e8aa0",-- -5974
x"d3a20",-- -11358
x"d46a0",-- -11158
x"db230",-- -9437
x"e0190",-- -8167
x"e6880",-- -6520
x"f17f0",-- -3713
x"f8070",-- -2041
x"f65c0",-- -2468
x"f5a70",-- -2649
x"f6ff0",-- -2305
x"f8a80",-- -1880
x"00980",-- 152
x"0eb10",-- 3761
x"1b4e0",-- 6990
x"1c320",-- 7218
x"133a0",-- 4922
x"08e10",-- 2273
x"fd8f0",-- -625
x"f4da0",-- -2854
x"f0620",-- -3998
x"f17a0",-- -3718
x"f3c40",-- -3132
x"f3bd0",-- -3139
x"f2490",-- -3511
x"eb880",-- -5240
x"e2690",-- -7575
x"dbb30",-- -9293
x"db360",-- -9418
x"de830",-- -8573
x"e41a0",-- -7142
x"ecb40",-- -4940
x"f6c30",-- -2365
x"fe5f0",-- -417
x"00960",-- 150
x"ff830",-- -125
x"fdd10",-- -559
x"fe020",-- -510
x"00760",-- 118
x"033a0",-- 826
x"053d0",-- 1341
x"04170",-- 1047
x"ff7c0",-- -132
x"fa4b0",-- -1461
x"f4dc0",-- -2852
x"f1d40",-- -3628
x"f0940",-- -3948
x"f17a0",-- -3718
x"f44e0",-- -2994
x"f7b20",-- -2126
x"fa170",-- -1513
x"fb180",-- -1256
x"f94d0",-- -1715
x"f6f80",-- -2312
x"f8bb0",-- -1861
x"fccf0",-- -817
x"02670",-- 615
x"06bd0",-- 1725
x"0acd0",-- 2765
x"0d790",-- 3449
x"0d6d0",-- 3437
x"0b4c0",-- 2892
x"07c70",-- 1991
x"05380",-- 1336
x"03d60",-- 982
x"03970",-- 919
x"04200",-- 1056
x"04110",-- 1041
x"02e60",-- 742
x"02890",-- 649
x"01c20",-- 450
x"03680",-- 872
x"05b00",-- 1456
x"08fc0",-- 2300
x"0e5f0",-- 3679
x"12780",-- 4728
x"15c30",-- 5571
x"18b90",-- 6329
x"1bb70",-- 7095
x"1d1c0",-- 7452
x"1ebf0",-- 7871
x"1fd80",-- 8152
x"211c0",-- 8476
x"23fd0",-- 9213
x"287c0",-- 10364
x"2b3f0",-- 11071
x"29be0",-- 10686
x"22220",-- 8738
x"13ab0",-- 5035
x"f9130",-- -1773
x"de010",-- -8703
x"d5020",-- -11006
x"d9180",-- -9960
x"e0330",-- -8141
x"e5ce0",-- -6706
x"f13b0",-- -3781
x"fcf70",-- -777
x"00990",-- 153
x"00250",-- 37
x"ffa30",-- -93
x"fc5f0",-- -929
x"fa5c0",-- -1444
x"00260",-- 38
x"0c630",-- 3171
x"13630",-- 4963
x"11240",-- 4388
x"0ade0",-- 2782
x"00690",-- 105
x"f4e60",-- -2842
x"ec990",-- -4967
x"ea230",-- -5597
x"eb810",-- -5247
x"ee470",-- -4537
x"f2030",-- -3581
x"f2800",-- -3456
x"eea00",-- -4448
x"e8f30",-- -5901
x"e57f0",-- -6785
x"e2c40",-- -7484
x"e1f20",-- -7694
x"e68a0",-- -6518
x"ef510",-- -4271
x"f9db0",-- -1573
x"01310",-- 305
x"026e0",-- 622
x"00250",-- 37
x"fd530",-- -685
x"fcb40",-- -844
x"fcff0",-- -769
x"fdc70",-- -569
x"fe8f0",-- -369
x"fe8e0",-- -370
x"fd810",-- -639
x"fb070",-- -1273
x"f79c0",-- -2148
x"f3b00",-- -3152
x"f0f30",-- -3853
x"efd30",-- -4141
x"f2f00",-- -3344
x"f8a30",-- -1885
x"fe660",-- -410
x"ff360",-- -202
x"fdbd0",-- -579
x"fe190",-- -487
x"fef70",-- -265
x"00700",-- 112
x"022b0",-- 555
x"059e0",-- 1438
x"09ea0",-- 2538
x"0c890",-- 3209
x"0cac0",-- 3244
x"0a3c0",-- 2620
x"05800",-- 1408
x"00a30",-- 163
x"fdbd0",-- -579
x"fd6f0",-- -657
x"fec80",-- -312
x"00df0",-- 223
x"03a10",-- 929
x"05f30",-- 1523
x"06e50",-- 1765
x"078a0",-- 1930
x"08660",-- 2150
x"0ac50",-- 2757
x"0dc20",-- 3522
x"110e0",-- 4366
x"14a20",-- 5282
x"176f0",-- 5999
x"19aa0",-- 6570
x"1bc80",-- 7112
x"1e270",-- 7719
x"1de10",-- 7649
x"1d9c0",-- 7580
x"1f000",-- 7936
x"240a0",-- 9226
x"27470",-- 10055
x"28040",-- 10244
x"24f10",-- 9457
x"192e0",-- 6446
x"00a00",-- 160
x"e46c0",-- -7060
x"d8230",-- -10205
x"d8640",-- -10140
x"da6e0",-- -9618
x"df900",-- -8304
x"f0c60",-- -3898
x"04910",-- 1169
x"0d5d0",-- 3421
x"0cd70",-- 3287
x"08fc0",-- 2300
x"00670",-- 103
x"f75b0",-- -2213
x"f80f0",-- -2033
x"00960",-- 150
x"06f90",-- 1785
x"08fe0",-- 2302
x"0a630",-- 2659
x"07650",-- 1893
x"fd340",-- -716
x"f0260",-- -4058
x"e65a0",-- -6566
x"e2d50",-- -7467
x"e4850",-- -7035
x"eb740",-- -5260
x"f3e50",-- -3099
x"f7b80",-- -2120
x"f5590",-- -2727
x"f0df0",-- -3873
x"eac10",-- -5439
x"e3e50",-- -7195
x"df720",-- -8334
x"e3b30",-- -7245
x"eeb10",-- -4431
x"f9fb0",-- -1541
x"01990",-- 409
x"05d10",-- 1489
x"063f0",-- 1599
x"03e70",-- 999
x"ff110",-- -239
x"fa3a0",-- -1478
x"f75e0",-- -2210
x"f7810",-- -2175
x"fa3f0",-- -1473
x"fcfc0",-- -772
x"fde00",-- -544
x"fb740",-- -1164
x"f7750",-- -2187
x"f2df0",-- -3361
x"f0a70",-- -3929
x"f1d60",-- -3626
x"f5db0",-- -2597
x"faf80",-- -1288
x"01ab0",-- 427
x"056d0",-- 1389
x"05400",-- 1344
x"04960",-- 1174
x"03ef0",-- 1007
x"03fe0",-- 1022
x"052e0",-- 1326
x"07060",-- 1798
x"098b0",-- 2443
x"0a900",-- 2704
x"08d70",-- 2263
x"05b20",-- 1458
x"00cb0",-- 203
x"fc910",-- -879
x"fa550",-- -1451
x"fb7e0",-- -1154
x"ff270",-- -217
x"03990",-- 921
x"07e00",-- 2016
x"0aef0",-- 2799
x"0d7c0",-- 3452
x"0d970",-- 3479
x"0cb10",-- 3249
x"0c540",-- 3156
x"0d990",-- 3481
x"116c0",-- 4460
x"16d70",-- 5847
x"19b90",-- 6585
x"1c2c0",-- 7212
x"1d7d0",-- 7549
x"1d290",-- 7465
x"1d960",-- 7574
x"1dab0",-- 7595
x"1ff80",-- 8184
x"21780",-- 8568
x"234e0",-- 9038
x"21dc0",-- 8668
x"17560",-- 5974
x"00640",-- 100
x"e8e60",-- -5914
x"de690",-- -8599
x"dd9f0",-- -8801
x"de560",-- -8618
x"e1000",-- -7936
x"ee5d0",-- -4515
x"025d0",-- 605
x"10570",-- 4183
x"11990",-- 4505
x"0b080",-- 2824
x"01180",-- 280
x"fb1a0",-- -1254
x"f9660",-- -1690
x"f9d00",-- -1584
x"fb7e0",-- -1154
x"ff290",-- -215
x"04a00",-- 1184
x"068c0",-- 1676
x"01fd0",-- 509
x"f65f0",-- -2465
x"ea320",-- -5582
x"e3fb0",-- -7173
x"e58e0",-- -6770
x"e98d0",-- -5747
x"ec8e0",-- -4978
x"ef100",-- -4336
x"f3930",-- -3181
x"f6a20",-- -2398
x"f2f50",-- -3339
x"ead70",-- -5417
x"e4100",-- -7152
x"e4b70",-- -6985
x"ea380",-- -5576
x"f2190",-- -3559
x"f9420",-- -1726
x"00530",-- 83
x"06660",-- 1638
x"0a460",-- 2630
x"08d10",-- 2257
x"01bd0",-- 445
x"fa110",-- -1519
x"f56f0",-- -2705
x"f54d0",-- -2739
x"f6be0",-- -2370
x"f7e70",-- -2073
x"f8350",-- -1995
x"f9cc0",-- -1588
x"faa00",-- -1376
x"f88a0",-- -1910
x"f59f0",-- -2657
x"f4550",-- -2987
x"f6d50",-- -2347
x"faf80",-- -1288
x"00000",-- 0
x"05760",-- 1398
x"09270",-- 2343
x"0ae50",-- 2789
x"0bf40",-- 3060
x"0b830",-- 2947
x"08db0",-- 2267
x"04340",-- 1076
x"00800",-- 128
x"ff6c0",-- -148
x"ff440",-- -188
x"fed70",-- -297
x"fe760",-- -394
x"ff2b0",-- -213
x"00b60",-- 182
x"01f60",-- 502
x"027a0",-- 634
x"03040",-- 772
x"04f20",-- 1266
x"084d0",-- 2125
x"0bf30",-- 3059
x"0e700",-- 3696
x"104a0",-- 4170
x"117e0",-- 4478
x"12520",-- 4690
x"133a0",-- 4922
x"13880",-- 5000
x"13870",-- 4999
x"14840",-- 5252
x"165e0",-- 5726
x"1a140",-- 6676
x"1df80",-- 7672
x"20460",-- 8262
x"22200",-- 8736
x"22e20",-- 8930
x"23530",-- 9043
x"20610",-- 8289
x"12c30",-- 4803
x"fac30",-- -1341
x"e7c00",-- -6208
x"e2670",-- -7577
x"e2c30",-- -7485
x"deab0",-- -8533
x"e17c0",-- -7812
x"f2d00",-- -3376
x"066e0",-- 1646
x"0f2c0",-- 3884
x"0e370",-- 3639
x"09fe0",-- 2558
x"03a40",-- 932
x"fcd20",-- -814
x"f7f30",-- -2061
x"f5bd0",-- -2627
x"f5ae0",-- -2642
x"fa480",-- -1464
x"01740",-- 372
x"05510",-- 1361
x"01740",-- 372
x"f8b10",-- -1871
x"f0e80",-- -3864
x"ebe50",-- -5147
x"e85d0",-- -6051
x"e5cf0",-- -6705
x"e58e0",-- -6770
x"e8de0",-- -5922
x"efe00",-- -4128
x"f4ee0",-- -2834
x"f3630",-- -3229
x"ee240",-- -4572
x"eae40",-- -5404
x"eb920",-- -5230
x"ece30",-- -4893
x"ee1e0",-- -4578
x"f2100",-- -3568
x"fb4d0",-- -1203
x"063e0",-- 1598
x"0ca50",-- 3237
x"0ba40",-- 2980
x"06ea0",-- 1770
x"01580",-- 344
x"fbe50",-- -1051
x"f5b10",-- -2639
x"f0c10",-- -3903
x"ee9b0",-- -4453
x"f09e0",-- -3938
x"f65c0",-- -2468
x"fb340",-- -1228
x"fc1e0",-- -994
x"fad20",-- -1326
x"fba90",-- -1111
x"fe730",-- -397
x"fe580",-- -424
x"fdb00",-- -592
x"00280",-- 40
x"05d10",-- 1489
x"0b130",-- 2835
x"0d180",-- 3352
x"0c570",-- 3159
x"09b00",-- 2480
x"04c80",-- 1224
x"00500",-- 80
x"fc6c0",-- -916
x"f9450",-- -1723
x"f8c60",-- -1850
x"fb9c0",-- -1124
x"00960",-- 150
x"05080",-- 1288
x"073a0",-- 1850
x"07bc0",-- 1980
x"08a70",-- 2215
x"08720",-- 2162
x"07ef0",-- 2031
x"066b0",-- 1643
x"065d0",-- 1629
x"08fe0",-- 2302
x"0ccf0",-- 3279
x"0eea0",-- 3818
x"104a0",-- 4170
x"12900",-- 4752
x"14dc0",-- 5340
x"15fd0",-- 5629
x"16570",-- 5719
x"17d20",-- 6098
x"1a250",-- 6693
x"1d880",-- 7560
x"1f290",-- 7977
x"205e0",-- 8286
x"21510",-- 8529
x"23190",-- 8985
x"1f580",-- 8024
x"0f990",-- 3993
x"fa850",-- -1403
x"ed1b0",-- -4837
x"e8530",-- -6061
x"e1970",-- -7785
x"db5a0",-- -9382
x"e1930",-- -7789
x"f3e30",-- -3101
x"03fb0",-- 1019
x"0b850",-- 2949
x"0e050",-- 3589
x"0d990",-- 3481
x"0a1b0",-- 2587
x"03f40",-- 1012
x"fb6d0",-- -1171
x"f3a70",-- -3161
x"f25f0",-- -3489
x"f7740",-- -2188
x"fd8a0",-- -630
x"ff800",-- -128
x"fe910",-- -367
x"fc3c0",-- -964
x"f81b0",-- -2021
x"f1e50",-- -3611
x"eb240",-- -5340
x"e5340",-- -6860
x"e2190",-- -7655
x"e4c60",-- -6970
x"eb700",-- -5264
x"ef4a0",-- -4278
x"ef400",-- -4288
x"f0320",-- -4046
x"f2dc0",-- -3364
x"f4080",-- -3064
x"f1480",-- -3768
x"efc90",-- -4151
x"f2eb0",-- -3349
x"fa3c0",-- -1476
x"01420",-- 322
x"054c0",-- 1356
x"06a20",-- 1698
x"07260",-- 1830
x"058f0",-- 1423
x"00350",-- 53
x"f93e0",-- -1730
x"f2800",-- -3456
x"ef520",-- -4270
x"f0060",-- -4090
x"f3200",-- -3296
x"f6320",-- -2510
x"f8fd0",-- -1795
x"fca70",-- -857
x"00260",-- 38
x"02080",-- 520
x"01360",-- 310
x"00de0",-- 222
x"02840",-- 644
x"05170",-- 1303
x"06cd0",-- 1741
x"07080",-- 1800
x"06b90",-- 1721
x"066e0",-- 1646
x"04db0",-- 1243
x"01c60",-- 454
x"fe730",-- -397
x"fc140",-- -1004
x"fc4d0",-- -947
x"fdb20",-- -590
x"ff800",-- -128
x"01bc0",-- 444
x"04780",-- 1144
x"06dc0",-- 1756
x"07c70",-- 1991
x"07310",-- 1841
x"062f0",-- 1583
x"06020",-- 1538
x"06570",-- 1623
x"07a90",-- 1961
x"09180",-- 2328
x"09ea0",-- 2538
x"0b2c0",-- 2860
x"0e8c0",-- 3724
x"12eb0",-- 4843
x"164f0",-- 5711
x"18500",-- 6224
x"1bb00",-- 7088
x"1f140",-- 7956
x"20e20",-- 8418
x"20370",-- 8247
x"1dc40",-- 7620
x"1c1b0",-- 7195
x"1bd00",-- 7120
x"1c400",-- 7232
x"15bf0",-- 5567
x"07040",-- 1796
x"f8e80",-- -1816
x"f2a80",-- -3416
x"ed7c0",-- -4740
x"e3130",-- -7405
x"dd410",-- -8895
x"e6cd0",-- -6451
x"f6e10",-- -2335
x"00a80",-- 168
x"05b30",-- 1459
x"0b590",-- 2905
x"0f6d0",-- 3949
x"0dec0",-- 3564
x"07170",-- 1815
x"fd2e0",-- -722
x"f5b50",-- -2635
x"f4e90",-- -2839
x"f7360",-- -2250
x"f7770",-- -2185
x"f6b60",-- -2378
x"f8e10",-- -1823
x"fba60",-- -1114
x"f9e20",-- -1566
x"f4410",-- -3007
x"eea70",-- -4441
x"ea550",-- -5547
x"e7560",-- -6314
x"e6aa0",-- -6486
x"e7920",-- -6254
x"e8240",-- -6108
x"e9f60",-- -5642
x"ee980",-- -4456
x"f37f0",-- -3201
x"f5430",-- -2749
x"f4de0",-- -2850
x"f6a80",-- -2392
x"fb180",-- -1256
x"fe9e0",-- -354
x"ff770",-- -137
x"fff60",-- -10
x"02160",-- 534
x"03c10",-- 961
x"01c40",-- 452
x"fd950",-- -619
x"f9cc0",-- -1588
x"f72f0",-- -2257
x"f5220",-- -2782
x"f39a0",-- -3174
x"f2c50",-- -3387
x"f3f30",-- -3085
x"f7240",-- -2268
x"fb250",-- -1243
x"fdd50",-- -555
x"00320",-- 50
x"02b40",-- 692
x"04a20",-- 1186
x"06280",-- 1576
x"067b0",-- 1659
x"05da0",-- 1498
x"048c0",-- 1164
x"03bd0",-- 957
x"03490",-- 841
x"01ec0",-- 492
x"00410",-- 65
x"ff170",-- -233
x"ff7b0",-- -133
x"00080",-- 8
x"003e0",-- 62
x"00840",-- 132
x"01ea0",-- 490
x"040c0",-- 1036
x"05010",-- 1281
x"04c70",-- 1223
x"04b10",-- 1201
x"05600",-- 1376
x"057c0",-- 1404
x"05440",-- 1348
x"054a0",-- 1354
x"069a0",-- 1690
x"08770",-- 2167
x"0a8e0",-- 2702
x"0d630",-- 3427
x"11210",-- 4385
x"149b0",-- 5275
x"17e40",-- 6116
x"1a0f0",-- 6671
x"1c140",-- 7188
x"1c610",-- 7265
x"1b9c0",-- 7068
x"1aa00",-- 6816
x"19300",-- 6448
x"19c90",-- 6601
x"1a9a0",-- 6810
x"1aed0",-- 6893
x"15bf0",-- 5567
x"0ab90",-- 2745
x"ff580",-- -168
x"f7180",-- -2280
x"ef790",-- -4231
x"e4f80",-- -6920
x"e04c0",-- -8116
x"e68c0",-- -6516
x"f2c30",-- -3389
x"facf0",-- -1329
x"00c10",-- 193
x"092c0",-- 2348
x"0f7e0",-- 3966
x"0f100",-- 3856
x"08190",-- 2073
x"00c80",-- 200
x"fbad0",-- -1107
x"f8820",-- -1918
x"f6000",-- -2560
x"f3d80",-- -3112
x"f3cf0",-- -3121
x"f6d00",-- -2352
x"f9ec0",-- -1556
x"f9110",-- -1775
x"f5520",-- -2734
x"f2cd0",-- -3379
x"f0ca0",-- -3894
x"ec380",-- -5064
x"e7400",-- -6336
x"e5a20",-- -6750
x"e6df0",-- -6433
x"e7e30",-- -6173
x"ea820",-- -5502
x"ef720",-- -4238
x"f4890",-- -2935
x"f7ea0",-- -2070
x"faa50",-- -1371
x"fe320",-- -462
x"003c0",-- 60
x"00660",-- 102
x"00030",-- 3
x"ffea0",-- -22
x"ff5d0",-- -163
x"fdf40",-- -524
x"fc3f0",-- -961
x"fa8e0",-- -1394
x"f8eb0",-- -1813
x"f7a90",-- -2135
x"f6520",-- -2478
x"f52a0",-- -2774
x"f5680",-- -2712
x"f73b0",-- -2245
x"f9510",-- -1711
x"fba40",-- -1116
x"fe620",-- -414
x"01c90",-- 457
x"04e30",-- 1251
x"07440",-- 1860
x"07c70",-- 1991
x"06300",-- 1584
x"05530",-- 1363
x"04200",-- 1056
x"01590",-- 345
x"fef30",-- -269
x"fe500",-- -432
x"feff0",-- -257
x"ffb20",-- -78
x"01270",-- 295
x"02f40",-- 756
x"043f0",-- 1087
x"05270",-- 1319
x"05950",-- 1429
x"04780",-- 1144
x"02710",-- 625
x"01270",-- 295
x"00a80",-- 168
x"00410",-- 65
x"003a0",-- 58
x"020f0",-- 527
x"05090",-- 1289
x"07ec0",-- 2028
x"0b1d0",-- 2845
x"0e7a0",-- 3706
x"11800",-- 4480
x"13e90",-- 5097
x"15fa0",-- 5626
x"179c0",-- 6044
x"17b50",-- 6069
x"17960",-- 6038
x"17850",-- 6021
x"17290",-- 5929
x"16980",-- 5784
x"16980",-- 5784
x"17170",-- 5911
x"17e70",-- 6119
x"19470",-- 6471
x"18e10",-- 6369
x"12040",-- 4612
x"073b0",-- 1851
x"fdcb0",-- -565
x"f8230",-- -2013
x"ef110",-- -4335
x"e4f10",-- -6927
x"e3b60",-- -7242
x"ec330",-- -5069
x"f5950",-- -2667
x"faaa0",-- -1366
x"01ab0",-- 427
x"0afe0",-- 2814
x"0f600",-- 3936
x"0d400",-- 3392
x"06dc0",-- 1756
x"ffd30",-- -45
x"fa1b0",-- -1509
x"f6700",-- -2448
x"f2c30",-- -3389
x"ee5f0",-- -4513
x"ef220",-- -4318
x"f4bb0",-- -2885
x"f83a0",-- -1990
x"f6c30",-- -2365
x"f6940",-- -2412
x"f8140",-- -2028
x"f6480",-- -2488
x"f0150",-- -4075
x"eacf0",-- -5425
x"e89b0",-- -5989
x"e7f90",-- -6151
x"e7110",-- -6383
x"e8260",-- -6106
x"ebfc0",-- -5124
x"f1fb0",-- -3589
x"f7e70",-- -2073
x"fb850",-- -1147
x"fecb0",-- -309
x"02030",-- 515
x"03d60",-- 982
x"026c0",-- 620
x"ff4e0",-- -178
x"fd160",-- -746
x"fb900",-- -1136
x"f9660",-- -1690
x"f7240",-- -2268
x"f6300",-- -2512
x"f6b10",-- -2383
x"f7f30",-- -2061
x"f8cf0",-- -1841
x"f9990",-- -1639
x"fad50",-- -1323
x"fd1b0",-- -741
x"febe0",-- -322
x"ff940",-- -108
x"00b70",-- 183
x"02ff0",-- 767
x"041c0",-- 1052
x"037c0",-- 892
x"03f30",-- 1011
x"045d0",-- 1117
x"03cc0",-- 972
x"02320",-- 562
x"018b0",-- 395
x"01590",-- 345
x"00b20",-- 178
x"00c30",-- 195
x"012c0",-- 300
x"01cc0",-- 460
x"027d0",-- 637
x"03760",-- 886
x"03dd0",-- 989
x"03590",-- 857
x"02db0",-- 731
x"027b0",-- 635
x"01bf0",-- 447
x"00c80",-- 200
x"01090",-- 265
x"02670",-- 615
x"04070",-- 1031
x"06640",-- 1636
x"09cb0",-- 2507
x"0d220",-- 3362
x"102f0",-- 4143
x"12a70",-- 4775
x"15180",-- 5400
x"16a20",-- 5794
x"16f40",-- 5876
x"15e60",-- 5606
x"14d60",-- 5334
x"13fb0",-- 5115
x"12410",-- 4673
x"112c0",-- 4396
x"11710",-- 4465
x"12870",-- 4743
x"14610",-- 5217
x"176c0",-- 5996
x"19320",-- 6450
x"15790",-- 5497
x"0d8a0",-- 3466
x"069f0",-- 1695
x"fff30",-- -13
x"f5ef0",-- -2577
x"ebfe0",-- -5122
x"e8800",-- -6016
x"ec0a0",-- -5110
x"f00d0",-- -4083
x"f4250",-- -3035
x"fa7a0",-- -1414
x"025c0",-- 604
x"07d30",-- 2003
x"08db0",-- 2267
x"06440",-- 1604
x"01fd0",-- 509
x"fe170",-- -489
x"fa020",-- -1534
x"f4460",-- -3002
x"ef4d0",-- -4275
x"eebb0",-- -4421
x"f1cc0",-- -3636
x"f3d90",-- -3111
x"f4a00",-- -2912
x"f7420",-- -2238
x"fa4b0",-- -1461
x"fa210",-- -1503
x"f5dd0",-- -2595
x"f0e10",-- -3871
x"ed150",-- -4843
x"e9dd0",-- -5667
x"e6fd0",-- -6403
x"e4e40",-- -6940
x"e68a0",-- -6518
x"ec0d0",-- -5107
x"f20a0",-- -3574
x"f73e0",-- -2242
x"fc700",-- -912
x"020a0",-- 522
x"05330",-- 1331
x"054f0",-- 1359
x"02ea0",-- 746
x"ff940",-- -108
x"fcaa0",-- -854
x"f9bf0",-- -1601
x"f6520",-- -2478
x"f3ed0",-- -3091
x"f4890",-- -2935
x"f7220",-- -2270
x"f9340",-- -1740
x"fb340",-- -1228
x"fe700",-- -400
x"01e00",-- 480
x"03670",-- 871
x"033d0",-- 829
x"027d0",-- 637
x"014a0",-- 330
x"000f0",-- 15
x"ff220",-- -222
x"fe690",-- -407
x"fe6e0",-- -402
x"feee0",-- -274
x"01490",-- 329
x"03680",-- 872
x"040f0",-- 1039
x"04750",-- 1141
x"05770",-- 1399
x"060f0",-- 1551
x"046c0",-- 1132
x"030b0",-- 779
x"027b0",-- 635
x"02120",-- 530
x"01150",-- 277
x"00440",-- 68
x"001e0",-- 30
x"00840",-- 132
x"01030",-- 259
x"01c60",-- 454
x"029b0",-- 667
x"03a80",-- 936
x"059f0",-- 1439
x"07db0",-- 2011
x"09ad0",-- 2477
x"0b360",-- 2870
x"0db70",-- 3511
x"0f920",-- 3986
x"10cd0",-- 4301
x"114f0",-- 4431
x"11fb0",-- 4603
x"124f0",-- 4687
x"11f80",-- 4600
x"11590",-- 4441
x"10550",-- 4181
x"10af0",-- 4271
x"11330",-- 4403
x"114c0",-- 4428
x"12c70",-- 4807
x"152b0",-- 5419
x"17e70",-- 6119
x"18c70",-- 6343
x"167c0",-- 5756
x"105a0",-- 4186
x"09770",-- 2423
x"03090",-- 777
x"f8be0",-- -1858
x"ee840",-- -4476
x"ea1c0",-- -5604
x"eada0",-- -5414
x"ec030",-- -5117
x"ee700",-- -4496
x"f58b0",-- -2677
x"fdc10",-- -575
x"03420",-- 834
x"06110",-- 1553
x"06aa0",-- 1706
x"05240",-- 1316
x"01740",-- 372
x"fcc80",-- -824
x"f7290",-- -2263
x"f1e50",-- -3611
x"ef970",-- -4201
x"efed0",-- -4115
x"f05d0",-- -4003
x"f1810",-- -3711
x"f5070",-- -2809
x"f8cf0",-- -1841
x"f99f0",-- -1633
x"f7a40",-- -2140
x"f50e0",-- -2802
x"f21e0",-- -3554
x"edd80",-- -4648
x"e8f70",-- -5897
x"e60d0",-- -6643
x"e6240",-- -6620
x"e84c0",-- -6068
x"ec230",-- -5085
x"f1ce0",-- -3634
x"f89e0",-- -1890
x"fee80",-- -280
x"04670",-- 1127
x"075b0",-- 1883
x"07180",-- 1816
x"052b0",-- 1323
x"02440",-- 580
x"fdb30",-- -589
x"f8800",-- -1920
x"f5340",-- -2764
x"f3e80",-- -3096
x"f3b30",-- -3149
x"f5650",-- -2715
x"f8e10",-- -1823
x"fcd40",-- -812
x"005c0",-- 92
x"035e0",-- 862
x"05150",-- 1301
x"05120",-- 1298
x"04230",-- 1059
x"024d0",-- 589
x"004e0",-- 78
x"feb20",-- -334
x"fe3e0",-- -450
x"fdfe0",-- -514
x"ff290",-- -215
x"02430",-- 579
x"04be0",-- 1214
x"06160",-- 1558
x"079e0",-- 1950
x"08a70",-- 2215
x"07df0",-- 2015
x"05b20",-- 1458
x"03da0",-- 986
x"01bf0",-- 447
x"ff7b0",-- -133
x"fe3a0",-- -454
x"fd720",-- -654
x"fde70",-- -537
x"ff220",-- -222
x"01670",-- 359
x"03850",-- 901
x"05970",-- 1431
x"079e0",-- 1950
x"09440",-- 2372
x"0a410",-- 2625
x"0a8b0",-- 2699
x"0af70",-- 2807
x"0b150",-- 2837
x"0b590",-- 2905
x"0ba40",-- 2980
x"0ca40",-- 3236
x"0ddd0",-- 3549
x"0f3a0",-- 3898
x"10130",-- 4115
x"10fa0",-- 4346
x"11f50",-- 4597
x"12270",-- 4647
x"125f0",-- 4703
x"12840",-- 4740
x"130d0",-- 4877
x"13240",-- 4900
x"14750",-- 5237
x"15c60",-- 5574
x"153b0",-- 5435
x"114a0",-- 4426
x"0c160",-- 3094
x"07dd0",-- 2013
x"01330",-- 307
x"f7a10",-- -2143
x"f03e0",-- -4034
x"ee2b0",-- -4565
x"ed270",-- -4825
x"eb630",-- -5277
x"ee4e0",-- -4530
x"f4980",-- -2920
x"fa3e0",-- -1474
x"fe2b0",-- -469
x"01c10",-- 449
x"03c90",-- 969
x"03150",-- 789
x"016c0",-- 364
x"fe580",-- -424
x"f97f0",-- -1665
x"f5590",-- -2727
x"f3930",-- -3181
x"f2530",-- -3501
x"f0750",-- -3979
x"f0960",-- -3946
x"f3470",-- -3257
x"f5040",-- -2812
x"f4a70",-- -2905
x"f3e50",-- -3099
x"f34a0",-- -3254
x"f1b30",-- -3661
x"eef00",-- -4368
x"ec4c0",-- -5044
x"eb1f0",-- -5345
x"ebfb0",-- -5125
x"ed520",-- -4782
x"ef5e0",-- -4258
x"f3cc0",-- -3124
x"f9750",-- -1675
x"fdd00",-- -560
x"01810",-- 385
x"046c0",-- 1132
x"04ef0",-- 1263
x"03da0",-- 986
x"01c90",-- 457
x"fe690",-- -407
x"fa170",-- -1513
x"f7750",-- -2187
x"f62f0",-- -2513
x"f5a90",-- -2647
x"f6840",-- -2428
x"f9510",-- -1711
x"fd270",-- -729
x"00320",-- 50
x"02940",-- 660
x"047f0",-- 1151
x"056c0",-- 1388
x"04ef0",-- 1263
x"03b80",-- 952
x"028e0",-- 654
x"01130",-- 275
x"00390",-- 57
x"00700",-- 112
x"018d0",-- 397
x"01e90",-- 489
x"03580",-- 856
x"05c40",-- 1476
x"06a50",-- 1701
x"05dd0",-- 1501
x"056f0",-- 1391
x"05b30",-- 1459
x"03ee0",-- 1006
x"01260",-- 294
x"001b0",-- 27
x"ff990",-- -103
x"fecb0",-- -309
x"fea50",-- -347
x"ffd30",-- -45
x"014a0",-- 330
x"02d10",-- 721
x"049d0",-- 1181
x"06300",-- 1584
x"07330",-- 1843
x"07fe0",-- 2046
x"08b30",-- 2227
x"08ef0",-- 2287
x"08ea0",-- 2282
x"09030",-- 2307
x"09b70",-- 2487
x"0a780",-- 2680
x"0b3b0",-- 2875
x"0c280",-- 3112
x"0d900",-- 3472
x"0eea0",-- 3818
x"0f920",-- 3986
x"104b0",-- 4171
x"11260",-- 4390
x"11a30",-- 4515
x"11eb0",-- 4587
x"12be0",-- 4798
x"13ec0",-- 5100
x"155a0",-- 5466
x"16630",-- 5731
x"15dd0",-- 5597
x"12220",-- 4642
x"0cb30",-- 3251
x"07800",-- 1920
x"002a0",-- 42
x"f6640",-- -2460
x"eeb40",-- -4428
x"ec780",-- -5000
x"ead70",-- -5417
x"e9720",-- -5774
x"eca00",-- -4960
x"f3950",-- -3179
x"f9560",-- -1706
x"fd580",-- -680
x"01d50",-- 469
x"04530",-- 1107
x"043c0",-- 1084
x"026e0",-- 622
x"ff4c0",-- -180
x"fa8e0",-- -1394
x"f62f0",-- -2513
x"f3650",-- -3227
x"f0f30",-- -3853
x"eef30",-- -4365
x"ef200",-- -4320
x"f19c0",-- -3684
x"f3ac0",-- -3156
x"f4980",-- -2920
x"f53b0",-- -2757
x"f6030",-- -2557
x"f56a0",-- -2710
x"f3380",-- -3272
x"f0780",-- -3976
x"eed70",-- -4393
x"ee350",-- -4555
x"ee0d0",-- -4595
x"ef160",-- -4330
x"f1a60",-- -3674
x"f5df0",-- -2593
x"fab20",-- -1358
x"ff090",-- -247
x"01d60",-- 470
x"03d30",-- 979
x"05630",-- 1379
x"04a00",-- 1184
x"01420",-- 322
x"fe0f0",-- -497
x"fc020",-- -1022
x"f98a0",-- -1654
x"f7330",-- -2253
x"f7100",-- -2288
x"f8690",-- -1943
x"faa30",-- -1373
x"fd880",-- -632
x"00750",-- 117
x"02bc0",-- 700
x"04fe0",-- 1278
x"06c20",-- 1730
x"06960",-- 1686
x"058f0",-- 1423
x"04b60",-- 1206
x"03df0",-- 991
x"02840",-- 644
x"01420",-- 322
x"01120",-- 274
x"01bd0",-- 445
x"02000",-- 512
x"02de0",-- 734
x"03f80",-- 1016
x"048f0",-- 1167
x"04700",-- 1136
x"04750",-- 1141
x"04620",-- 1122
x"02e00",-- 736
x"019a0",-- 410
x"014e0",-- 334
x"008f0",-- 143
x"ff6d0",-- -147
x"ff330",-- -205
x"00350",-- 53
x"00f40",-- 244
x"018a0",-- 394
x"033a0",-- 826
x"04e80",-- 1256
x"05f80",-- 1528
x"06fe0",-- 1790
x"081b0",-- 2075
x"08610",-- 2145
x"08a00",-- 2208
x"09510",-- 2385
x"09bc0",-- 2492
x"09ea0",-- 2538
x"0a960",-- 2710
x"0bd00",-- 3024
x"0cb80",-- 3256
x"0d7c0",-- 3452
x"0e0c0",-- 3596
x"0f380",-- 3896
x"102d0",-- 4141
x"10b80",-- 4280
x"11490",-- 4425
x"126b0",-- 4715
x"13c10",-- 5057
x"14db0",-- 5339
x"15970",-- 5527
x"143c0",-- 5180
x"10c30",-- 4291
x"0c1e0",-- 3102
x"076d0",-- 1901
x"fff80",-- -8
x"f75e0",-- -2210
x"f11d0",-- -3811
x"ee700",-- -4496
x"ec0f0",-- -5105
x"ea050",-- -5627
x"ecde0",-- -4898
x"f1ab0",-- -3669
x"f5720",-- -2702
x"f9450",-- -1723
x"fddb0",-- -549
x"004e0",-- 78
x"00d40",-- 212
x"01800",-- 384
x"00490",-- 73
x"fc500",-- -944
x"f91d0",-- -1763
x"f7590",-- -2215
x"f44e0",-- -2994
x"f1390",-- -3783
x"f0d70",-- -3881
x"f2610",-- -3487
x"f3110",-- -3311
x"f3900",-- -3184
x"f5330",-- -2765
x"f6690",-- -2455
x"f6340",-- -2508
x"f5380",-- -2760
x"f4170",-- -3049
x"f26c0",-- -3476
x"f12c0",-- -3796
x"f07a0",-- -3974
x"f0af0",-- -3921
x"f1ed0",-- -3603
x"f41e0",-- -3042
x"f6eb0",-- -2325
x"fa850",-- -1403
x"fe110",-- -495
x"008a0",-- 138
x"02ca0",-- 714
x"04710",-- 1137
x"03f10",-- 1009
x"021b0",-- 539
x"00ed0",-- 237
x"fead0",-- -339
x"fba30",-- -1117
x"f9fd0",-- -1539
x"f9830",-- -1661
x"f9150",-- -1771
x"f9d50",-- -1579
x"fbdb0",-- -1061
x"fdf10",-- -527
x"007a0",-- 122
x"03060",-- 774
x"052b0",-- 1323
x"068c0",-- 1676
x"077c0",-- 1916
x"07c20",-- 1986
x"07770",-- 1911
x"06b60",-- 1718
x"05740",-- 1396
x"042a0",-- 1066
x"03150",-- 789
x"02520",-- 594
x"01880",-- 392
x"011f0",-- 287
x"01d30",-- 467
x"01770",-- 375
x"00940",-- 148
x"01360",-- 310
x"015b0",-- 347
x"00410",-- 65
x"ffb80",-- -72
x"00840",-- 132
x"00080",-- 8
x"ff510",-- -175
x"003c0",-- 60
x"00cf0",-- 207
x"012c0",-- 300
x"02160",-- 534
x"033b0",-- 827
x"03f60",-- 1014
x"04f00",-- 1264
x"065a0",-- 1626
x"075d0",-- 1885
x"07f90",-- 2041
x"08b80",-- 2232
x"099a0",-- 2458
x"09f30",-- 2547
x"0a0a0",-- 2570
x"0a500",-- 2640
x"0b0e0",-- 2830
x"0b800",-- 2944
x"0b8b0",-- 2955
x"0c140",-- 3092
x"0cf90",-- 3321
x"0e130",-- 3603
x"0ef70",-- 3831
x"106b0",-- 4203
x"12c00",-- 4800
x"149a0",-- 5274
x"16340",-- 5684
x"169f0",-- 5791
x"14900",-- 5264
x"104f0",-- 4175
x"0bbc0",-- 3004
x"05560",-- 1366
x"fc2d0",-- -979
x"f42d0",-- -3027
x"ef3b0",-- -4293
x"eb2f0",-- -5329
x"e7830",-- -6269
x"e7bd0",-- -6211
x"eb700",-- -5264
x"ef6f0",-- -4241
x"f3ef0",-- -3089
x"f9200",-- -1760
x"fdf10",-- -527
x"01360",-- 310
x"03170",-- 791
x"036a0",-- 874
x"01cc0",-- 460
x"ff0b0",-- -245
x"fc2d0",-- -979
x"f8de0",-- -1826
x"f57e0",-- -2690
x"f2f80",-- -3336
x"f2490",-- -3511
x"f2ac0",-- -3412
x"f2e80",-- -3352
x"f37a0",-- -3206
x"f4cd0",-- -2867
x"f6140",-- -2540
x"f5f90",-- -2567
x"f5160",-- -2794
x"f4440",-- -3004
x"f3590",-- -3239
x"f1b30",-- -3661
x"f0a20",-- -3934
x"f11a0",-- -3814
x"f2350",-- -3531
x"f4260",-- -3034
x"f7f60",-- -2058
x"fbf30",-- -1037
x"ff040",-- -252
x"019e0",-- 414
x"04e60",-- 1254
x"06340",-- 1588
x"04d40",-- 1236
x"033d0",-- 829
x"01d00",-- 464
x"ff540",-- -172
x"fb8f0",-- -1137
x"f9770",-- -1673
x"f8ee0",-- -1810
x"f8410",-- -1983
x"f8d70",-- -1833
x"fabc0",-- -1348
x"fda30",-- -605
x"006b0",-- 107
x"04070",-- 1031
x"074a0",-- 1866
x"09330",-- 2355
x"0a590",-- 2649
x"0b0d0",-- 2829
x"0ab80",-- 2744
x"08c20",-- 2242
x"069f0",-- 1695
x"04ae0",-- 1198
x"02e00",-- 736
x"00660",-- 102
x"ff350",-- -203
x"fe620",-- -414
x"fe500",-- -432
x"fed50",-- -299
x"ff6d0",-- -147
x"fff30",-- -13
x"00800",-- 128
x"01770",-- 375
x"01720",-- 370
x"00f40",-- 244
x"00af0",-- 175
x"00b70",-- 183
x"003c0",-- 60
x"ffec0",-- -20
x"00200",-- 32
x"00fc0",-- 252
x"01bc0",-- 444
x"02940",-- 660
x"04190",-- 1049
x"051d0",-- 1309
x"061e0",-- 1566
x"07380",-- 1848
x"07c60",-- 1990
x"08000",-- 2048
x"087a0",-- 2170
x"08c00",-- 2240
x"088e0",-- 2190
x"08b40",-- 2228
x"09080",-- 2312
x"097e0",-- 2430
x"0a5f0",-- 2655
x"0b330",-- 2867
x"0c9f0",-- 3231
x"0e6d0",-- 3693
x"10a70",-- 4263
x"129a0",-- 4762
x"14e00",-- 5344
x"175a0",-- 5978
x"17c80",-- 6088
x"17060",-- 5894
x"132e0",-- 4910
x"0ee00",-- 3808
x"08ed0",-- 2285
x"005a0",-- 90
x"f7840",-- -2172
x"f0fa0",-- -3846
x"ecd90",-- -4903
x"e79d0",-- -6243
x"e5e30",-- -6685
x"e8c60",-- -5946
x"ec650",-- -5019
x"efd90",-- -4135
x"f5a20",-- -2654
x"fc070",-- -1017
x"fffe0",-- -2
x"02e60",-- 742
x"05630",-- 1379
x"05600",-- 1376
x"02980",-- 664
x"008f0",-- 143
x"fddb0",-- -549
x"f97a0",-- -1670
x"f5b80",-- -2632
x"f47d0",-- -2947
x"f3ac0",-- -3156
x"f2780",-- -3464
x"f2df0",-- -3361
x"f44b0",-- -2997
x"f5950",-- -2667
x"f6280",-- -2520
x"f6930",-- -2413
x"f65a0",-- -2470
x"f63e0",-- -2498
x"f5770",-- -2697
x"f4320",-- -3022
x"f36a0",-- -3222
x"f3bd0",-- -3139
x"f47b0",-- -2949
x"f5fb0",-- -2565
x"f8aa0",-- -1878
x"fb620",-- -1182
x"fe710",-- -399
x"01a40",-- 420
x"042a0",-- 1066
x"050b0",-- 1291
x"04e80",-- 1256
x"04820",-- 1154
x"02f20",-- 754
x"00140",-- 20
x"fd2f0",-- -721
x"fb450",-- -1211
x"f9e90",-- -1559
x"f85d0",-- -1955
x"f8a50",-- -1883
x"fa6c0",-- -1428
x"fca50",-- -859
x"ffb50",-- -75
x"03300",-- 816
x"068c0",-- 1676
x"08e10",-- 2273
x"0b010",-- 2817
x"0c000",-- 3072
x"0b720",-- 2930
x"09dd0",-- 2525
x"07d60",-- 2006
x"05830",-- 1411
x"029d0",-- 669
x"ffe90",-- -23
x"fdee0",-- -530
x"fd160",-- -746
x"fc930",-- -877
x"fcbe0",-- -834
x"fdc10",-- -575
x"ff300",-- -208
x"00940",-- 148
x"01830",-- 387
x"02390",-- 569
x"01b00",-- 432
x"00af0",-- 175
x"00230",-- 35
x"ff1f0",-- -225
x"fdef0",-- -529
x"fdcb0",-- -565
x"ff070",-- -249
x"fffb0",-- -5
x"00be0",-- 190
x"03100",-- 784
x"04f90",-- 1273
x"05f30",-- 1523
x"070b0",-- 1803
x"07c10",-- 1985
x"07ae0",-- 1966
x"07560",-- 1878
x"07030",-- 1795
x"068c0",-- 1676
x"06230",-- 1571
x"06210",-- 1569
x"06a90",-- 1705
x"079a0",-- 1946
x"08ff0",-- 2303
x"0ab30",-- 2739
x"0d090",-- 3337
x"0f2c0",-- 3884
x"118a0",-- 4490
x"13770",-- 4983
x"15d50",-- 5589
x"178f0",-- 6031
x"17a30",-- 6051
x"16ca0",-- 5834
x"13830",-- 4995
x"0f060",-- 3846
x"09180",-- 2328
x"02260",-- 550
x"f9cb0",-- -1589
x"f2c30",-- -3389
x"ee910",-- -4463
x"ea0b0",-- -5621
x"e6d80",-- -6440
x"e8120",-- -6126
x"eb7c0",-- -5252
x"ee240",-- -4572
x"f27d0",-- -3459
x"f85a0",-- -1958
x"fd240",-- -732
x"fffe0",-- -2
x"03560",-- 854
x"05040",-- 1284
x"03e70",-- 999
x"02c00",-- 704
x"017b0",-- 379
x"fe990",-- -359
x"fb100",-- -1264
x"f9b80",-- -1608
x"f88f0",-- -1905
x"f6bc0",-- -2372
x"f5d00",-- -2608
x"f62a0",-- -2518
x"f6190",-- -2535
x"f5c00",-- -2624
x"f5ac0",-- -2644
x"f4fd0",-- -2819
x"f4800",-- -2944
x"f3e50",-- -3099
x"f3360",-- -3274
x"f2910",-- -3439
x"f3110",-- -3311
x"f4170",-- -3049
x"f5c40",-- -2620
x"f83a0",-- -1990
x"fb2c0",-- -1236
x"fe960",-- -362
x"01f30",-- 499
x"05080",-- 1288
x"06cc0",-- 1740
x"08110",-- 2065
x"087a0",-- 2170
x"07810",-- 1921
x"04ca0",-- 1226
x"01c60",-- 454
x"fe430",-- -445
x"fb520",-- -1198
x"f7f40",-- -2060
x"f57e0",-- -2690
x"f5b50",-- -2635
x"f7480",-- -2232
x"f99f0",-- -1633
x"fc430",-- -957
x"018f0",-- 399
x"06140",-- 1556
x"08f20",-- 2290
x"0bba0",-- 3002
x"0d720",-- 3442
x"0ccf0",-- 3279
x"0b310",-- 2865
x"092b0",-- 2347
x"05860",-- 1414
x"017c0",-- 380
x"fec80",-- -312
x"fce60",-- -794
x"fa5a0",-- -1446
x"f9330",-- -1741
x"fa320",-- -1486
x"fb2c0",-- -1236
x"fbd10",-- -1071
x"fd7c0",-- -644
x"ff470",-- -185
x"00370",-- 55
x"00aa0",-- 170
x"00ed0",-- 237
x"00b70",-- 183
x"00200",-- 32
x"000f0",-- 15
x"ff650",-- -155
x"ff850",-- -123
x"00020",-- 2
x"00aa0",-- 170
x"01ef0",-- 495
x"03010",-- 769
x"04410",-- 1089
x"05ab0",-- 1451
x"06cd0",-- 1741
x"06f40",-- 1780
x"07a40",-- 1956
x"07e70",-- 2023
x"07a60",-- 1958
x"078f0",-- 1935
x"084d0",-- 2125
x"08aa0",-- 2218
x"09330",-- 2355
x"0a9f0",-- 2719
x"0c2a0",-- 3114
x"0e050",-- 3589
x"0fba0",-- 4026
x"11f00",-- 4592
x"14720",-- 5234
x"16cd0",-- 5837
x"17bf0",-- 6079
x"171c0",-- 5916
x"14950",-- 5269
x"11650",-- 4453
x"0c2d0",-- 3117
x"042f0",-- 1071
x"fc430",-- -957
x"f6000",-- -2560
x"f0660",-- -3994
x"ea080",-- -5624
x"e7220",-- -6366
x"e7470",-- -6329
x"e81f0",-- -6113
x"eaa50",-- -5467
x"ef020",-- -4350
x"f40c0",-- -3060
x"f8610",-- -1951
x"fd6f0",-- -657
x"01f10",-- 497
x"03f80",-- 1016
x"04aa0",-- 1194
x"060f0",-- 1551
x"05ab0",-- 1451
x"02ca0",-- 714
x"00440",-- 68
x"fef20",-- -270
x"fcbb0",-- -837
x"f9b70",-- -1609
x"f7df0",-- -2081
x"f6c50",-- -2363
x"f5980",-- -2664
x"f4670",-- -2969
x"f3ba0",-- -3142
x"f34a0",-- -3254
x"f2ff0",-- -3329
x"f2ad0",-- -3411
x"f2ad0",-- -3411
x"f2da0",-- -3366
x"f3200",-- -3296
x"f4500",-- -2992
x"f61c0",-- -2532
x"f7bf0",-- -2113
x"f9d80",-- -1576
x"fcee0",-- -786
x"ffdb0",-- -37
x"01f90",-- 505
x"04230",-- 1059
x"06190",-- 1561
x"06e10",-- 1761
x"07030",-- 1795
x"06bb0",-- 1723
x"05860",-- 1414
x"03ce0",-- 974
x"025d0",-- 605
x"00b10",-- 177
x"fda40",-- -604
x"fb9e0",-- -1122
x"fb390",-- -1223
x"fab60",-- -1354
x"f9e90",-- -1559
x"fb3e0",-- -1218
x"fe7f0",-- -385
x"00700",-- 112
x"026e0",-- 622
x"05530",-- 1363
x"071f0",-- 1823
x"07940",-- 1940
x"07d80",-- 2008
x"07220",-- 1826
x"04e10",-- 1249
x"030d0",-- 781
x"01a40",-- 420
x"ff9f0",-- -97
x"fd710",-- -655
x"fce30",-- -797
x"fcfa0",-- -774
x"fc9d0",-- -867
x"fca70",-- -857
x"fda10",-- -607
x"fecb0",-- -309
x"ff2b0",-- -213
x"ff8b0",-- -117
x"ffc90",-- -55
x"ffe00",-- -32
x"ff5d0",-- -163
x"fe340",-- -460
x"fdcc0",-- -564
x"fd940",-- -620
x"fd340",-- -716
x"fd7b0",-- -645
x"fec50",-- -315
x"002f0",-- 47
x"01740",-- 372
x"03ae0",-- 942
x"054c0",-- 1356
x"06440",-- 1604
x"07590",-- 1881
x"07ec0",-- 2028
x"078d0",-- 1933
x"07300",-- 1840
x"070b0",-- 1803
x"06c20",-- 1730
x"06cc0",-- 1740
x"07630",-- 1891
x"085a0",-- 2138
x"09b00",-- 2480
x"0bb20",-- 2994
x"0e000",-- 3584
x"109f0",-- 4255
x"13470",-- 4935
x"16700",-- 5744
x"18cc0",-- 6348
x"19be0",-- 6590
x"17f60",-- 6134
x"157d0",-- 5501
x"11f80",-- 4600
x"0b080",-- 2824
x"02d90",-- 729
x"fafc0",-- -1284
x"f5740",-- -2700
x"ee2b0",-- -4565
x"e88d0",-- -6003
x"e6300",-- -6608
x"e5e50",-- -6683
x"e6fc0",-- -6404
x"e9720",-- -5774
x"edcc0",-- -4660
x"f1ed0",-- -3603
x"f76f0",-- -2193
x"fc750",-- -907
x"00020",-- 2
x"02430",-- 579
x"05120",-- 1298
x"06a20",-- 1698
x"05e90",-- 1513
x"04a50",-- 1189
x"03a10",-- 929
x"02d40",-- 724
x"006b0",-- 107
x"fe5c0",-- -420
x"fc4d0",-- -947
x"fad90",-- -1319
x"f8e90",-- -1815
x"f6f70",-- -2313
x"f5100",-- -2800
x"f3a40",-- -3164
x"f2930",-- -3437
x"f1560",-- -3754
x"f0bb0",-- -3909
x"f0370",-- -4041
x"f0f30",-- -3853
x"f20a0",-- -3574
x"f3f60",-- -3082
x"f5b80",-- -2632
x"f8940",-- -1900
x"fbd00",-- -1072
x"fee60",-- -282
x"01620",-- 354
x"038d0",-- 909
x"05b00",-- 1456
x"06e30",-- 1763
x"078d0",-- 1933
x"07670",-- 1895
x"06f90",-- 1785
x"063e0",-- 1598
x"05a90",-- 1449
x"04b10",-- 1201
x"03630",-- 867
x"02490",-- 585
x"01720",-- 370
x"00c50",-- 197
x"00000",-- 0
x"ff2c0",-- -212
x"feb90",-- -327
x"fecf0",-- -305
x"fed70",-- -297
x"fea30",-- -349
x"feac0",-- -340
x"ff420",-- -190
x"ff7c0",-- -132
x"ff9c0",-- -100
x"ff860",-- -122
x"ff6a0",-- -150
x"ffb20",-- -78
x"000f0",-- 15
x"00350",-- 53
x"001e0",-- 30
x"00af0",-- 175
x"013b0",-- 315
x"017e0",-- 382
x"01220",-- 290
x"01100",-- 272
x"00700",-- 112
x"ff830",-- -125
x"fe8f0",-- -369
x"fd3d0",-- -707
x"fc1c0",-- -996
x"fb5b0",-- -1189
x"fb5b0",-- -1189
x"fb020",-- -1278
x"fb4f0",-- -1201
x"fc5f0",-- -929
x"fd9a0",-- -614
x"fefc0",-- -260
x"00840",-- 132
x"01f10",-- 497
x"03380",-- 824
x"04760",-- 1142
x"05090",-- 1289
x"05670",-- 1383
x"05790",-- 1401
x"05970",-- 1431
x"05920",-- 1426
x"05970",-- 1431
x"05d50",-- 1493
x"069f0",-- 1695
x"082b0",-- 2091
x"09a10",-- 2465
x"0b920",-- 2962
x"0dd50",-- 3541
x"10870",-- 4231
x"13240",-- 4900
x"15d00",-- 5584
x"18890",-- 6281
x"1aae0",-- 6830
x"1b1c0",-- 6940
x"19260",-- 6438
x"165e0",-- 5726
x"12640",-- 4708
x"0bab0",-- 2987
x"03600",-- 864
x"fc930",-- -877
x"f6a80",-- -2392
x"ef7c0",-- -4228
x"ea170",-- -5609
x"e7d60",-- -6186
x"e6d00",-- -6448
x"e6670",-- -6553
x"e8600",-- -6048
x"eb7a0",-- -5254
x"ee9b0",-- -4453
x"f31f0",-- -3297
x"f7d50",-- -2091
x"fb720",-- -1166
x"fec50",-- -315
x"02ac0",-- 684
x"051d0",-- 1309
x"060d0",-- 1549
x"06e00",-- 1760
x"07a60",-- 1958
x"07310",-- 1841
x"05c10",-- 1473
x"04440",-- 1092
x"02460",-- 582
x"ffbf0",-- -65
x"fca20",-- -862
x"f9c60",-- -1594
x"f6c50",-- -2363
x"f3e50",-- -3099
x"f14c0",-- -3764
x"ef630",-- -4253
x"ee4e0",-- -4530
x"ed880",-- -4728
x"edb60",-- -4682
x"ef130",-- -4333
x"f0fc0",-- -3844
x"f2e30",-- -3357
x"f5b30",-- -2637
x"f8df0",-- -1825
x"fb920",-- -1134
x"fe440",-- -444
x"00cb0",-- 203
x"02f00",-- 752
x"04bb0",-- 1211
x"06780",-- 1656
x"07630",-- 1891
x"08210",-- 2081
x"08ed0",-- 2285
x"09510",-- 2385
x"09330",-- 2355
x"08e60",-- 2278
x"08c00",-- 2240
x"072c0",-- 1836
x"05680",-- 1384
x"042d0",-- 1069
x"01a90",-- 425
x"fea80",-- -344
x"fcde0",-- -802
x"fc730",-- -909
x"fa370",-- -1481
x"f9450",-- -1723
x"f9e50",-- -1563
x"fa110",-- -1519
x"fa840",-- -1404
x"fb850",-- -1147
x"fca00",-- -864
x"fd710",-- -655
x"ff490",-- -183
x"003a0",-- 58
x"00f20",-- 242
x"01cc0",-- 460
x"02f00",-- 752
x"03530",-- 851
x"02d70",-- 727
x"02750",-- 629
x"022b0",-- 555
x"01a80",-- 424
x"006b0",-- 107
x"ff860",-- -122
x"febe0",-- -322
x"fe390",-- -455
x"fdb20",-- -590
x"fd160",-- -746
x"fca50",-- -859
x"fcad0",-- -851
x"fcd40",-- -812
x"fd2f0",-- -721
x"fdd50",-- -555
x"fe490",-- -439
x"ff880",-- -120
x"00ad0",-- 173
x"018a0",-- 394
x"020a0",-- 522
x"032e0",-- 814
x"040a0",-- 1034
x"04c20",-- 1218
x"05920",-- 1426
x"06440",-- 1604
x"07ae0",-- 1966
x"09440",-- 2372
x"0ad40",-- 2772
x"0ca20",-- 3234
x"0ef40",-- 3828
x"11360",-- 4406
x"13a10",-- 5025
x"160c0",-- 5644
x"18540",-- 6228
x"19fb0",-- 6651
x"1aac0",-- 6828
x"19040",-- 6404
x"16a50",-- 5797
x"12d40",-- 4820
x"0cdc0",-- 3292
x"05e70",-- 1511
x"ff670",-- -153
x"f9600",-- -1696
x"f2460",-- -3514
x"ed400",-- -4800
x"e9a60",-- -5722
x"e78e0",-- -6258
x"e6330",-- -6605
x"e6e90",-- -6423
x"e8aa0",-- -5974
x"eb040",-- -5372
x"eed70",-- -4393
x"f2af0",-- -3409
x"f6b60",-- -2378
x"fa640",-- -1436
x"fea00",-- -352
x"018b0",-- 395
x"03ea0",-- 1002
x"05ea0",-- 1514
x"07620",-- 1890
x"07f80",-- 2040
x"07a90",-- 1961
x"07490",-- 1865
x"05c90",-- 1481
x"04140",-- 1044
x"01a30",-- 419
x"ff400",-- -192
x"fc5a0",-- -934
x"f9630",-- -1693
x"f6890",-- -2423
x"f41e0",-- -3042
x"f2250",-- -3547
x"f03f0",-- -4033
x"ef570",-- -4265
x"eefa0",-- -4358
x"ef480",-- -4280
x"efb80",-- -4168
x"f1400",-- -3776
x"f3010",-- -3327
x"f5240",-- -2780
x"f78d0",-- -2163
x"fa140",-- -1516
x"fcc60",-- -826
x"ff6d0",-- -147
x"02460",-- 582
x"04a90",-- 1193
x"07220",-- 1826
x"09490",-- 2377
x"0b1a0",-- 2842
x"0c450",-- 3141
x"0d2e0",-- 3374
x"0d8b0",-- 3467
x"0cca0",-- 3274
x"0b990",-- 2969
x"09800",-- 2432
x"06500",-- 1616
x"034c0",-- 844
x"00eb0",-- 235
x"fe390",-- -455
x"fb1a0",-- -1254
x"fa110",-- -1519
x"f94f0",-- -1713
x"f8760",-- -1930
x"f8140",-- -2028
x"f8610",-- -1951
x"f92e0",-- -1746
x"f9cb0",-- -1589
x"fad50",-- -1323
x"fb740",-- -1164
x"fccf0",-- -817
x"fe460",-- -442
x"ff9a0",-- -102
x"00b60",-- 182
x"01670",-- 359
x"02870",-- 647
x"031a0",-- 794
x"03470",-- 839
x"03240",-- 804
x"032c0",-- 812
x"02b40",-- 692
x"020a0",-- 522
x"01290",-- 297
x"00230",-- 35
x"ff740",-- -140
x"feb40",-- -332
x"fe640",-- -412
x"fe2b0",-- -469
x"fe300",-- -464
x"fe3a0",-- -454
x"ff360",-- -202
x"ffd80",-- -40
x"00760",-- 118
x"01710",-- 369
x"02890",-- 649
x"036c0",-- 876
x"044d0",-- 1101
x"054a0",-- 1354
x"06500",-- 1616
x"07f30",-- 2035
x"09740",-- 2420
x"0b2c0",-- 2860
x"0d580",-- 3416
x"0fc40",-- 4036
x"12870",-- 4743
x"15730",-- 5491
x"185a0",-- 6234
x"1ad70",-- 6871
x"1c630",-- 7267
x"1ba80",-- 7080
x"1a130",-- 6675
x"17600",-- 5984
x"12110",-- 4625
x"0b880",-- 2952
x"05120",-- 1298
x"ff1a0",-- -230
x"f7e70",-- -2073
x"f1ed0",-- -3603
x"ecbc0",-- -4932
x"ea850",-- -5499
x"e7160",-- -6378
x"e6920",-- -6510
x"e7a60",-- -6234
x"e8320",-- -6094
x"eb240",-- -5340
x"ee100",-- -4592
x"f0fc0",-- -3844
x"f4bc0",-- -2884
x"f88a0",-- -1910
x"fb7e0",-- -1154
x"feac0",-- -340
x"006e0",-- 110
x"03850",-- 901
x"04850",-- 1157
x"06070",-- 1543
x"06e10",-- 1761
x"06a50",-- 1701
x"06e50",-- 1765
x"05950",-- 1429
x"04ed0",-- 1261
x"034f0",-- 847
x"00e10",-- 225
x"fe820",-- -382
x"fbf60",-- -1034
x"f99a0",-- -1638
x"f6700",-- -2448
x"f41b0",-- -3045
x"f26c0",-- -3476
x"f0c50",-- -3899
x"efae0",-- -4178
x"eefc0",-- -4356
x"ef3b0",-- -4293
x"f0290",-- -4055
x"f1290",-- -3799
x"f2fd0",-- -3331
x"f4fc0",-- -2820
x"f7650",-- -2203
x"fa3f0",-- -1473
x"fd310",-- -719
x"00390",-- 57
x"03090",-- 777
x"062d0",-- 1581
x"08d70",-- 2263
x"0b470",-- 2887
x"0cff0",-- 3327
x"0d8a0",-- 3466
x"0d630",-- 3427
x"0caf0",-- 3247
x"0b920",-- 2962
x"09290",-- 2345
x"070e0",-- 1806
x"052e0",-- 1326
x"03670",-- 871
x"014c0",-- 332
x"ff440",-- -188
x"fdea0",-- -534
x"fc7a0",-- -902
x"fb470",-- -1209
x"fa0f0",-- -1521
x"f9480",-- -1720
x"f8a80",-- -1880
x"f87a0",-- -1926
x"f8cd0",-- -1843
x"f9610",-- -1695
x"fa4e0",-- -1458
x"fb900",-- -1136
x"fd060",-- -762
x"fe800",-- -384
x"ffe70",-- -25
x"011c0",-- 284
x"024b0",-- 587
x"03150",-- 789
x"03ab0",-- 939
x"03cc0",-- 972
x"036f0",-- 879
x"02d40",-- 724
x"02670",-- 615
x"01df0",-- 479
x"010d0",-- 269
x"00870",-- 135
x"00850",-- 133
x"00940",-- 148
x"00c50",-- 197
x"010b0",-- 267
x"01810",-- 385
x"020a0",-- 522
x"02690",-- 617
x"02c80",-- 712
x"02c80",-- 712
x"03300",-- 816
x"03b70",-- 951
x"04a20",-- 1186
x"05a80",-- 1448
x"06f40",-- 1780
x"08e80",-- 2280
x"0b2c0",-- 2860
x"0ddd0",-- 3549
x"10ae0",-- 4270
x"13b00",-- 5040
x"16660",-- 5734
x"18a20",-- 6306
x"197d0",-- 6525
x"191a0",-- 6426
x"17cd0",-- 6093
x"14ef0",-- 5359
x"109a0",-- 4250
x"0b5b0",-- 2907
x"06550",-- 1621
x"00de0",-- 222
x"fb400",-- -1216
x"f62a0",-- -2518
x"f28f0",-- -3441
x"ef7e0",-- -4226
x"eccd0",-- -4915
x"eb4c0",-- -5300
x"eaac0",-- -5460
x"eb1a0",-- -5350
x"ebac0",-- -5204
x"ecd20",-- -4910
x"ee710",-- -4495
x"f0980",-- -3944
x"f2a50",-- -3419
x"f4b40",-- -2892
x"f6fa0",-- -2310
x"f94f0",-- -1713
x"fba90",-- -1111
x"fde00",-- -544
x"00120",-- 18
x"02030",-- 515
x"03b20",-- 946
x"04f90",-- 1273
x"05fe0",-- 1534
x"065a0",-- 1626
x"06210",-- 1569
x"05530",-- 1363
x"03f80",-- 1016
x"02340",-- 564
x"00000",-- 0
x"fd680",-- -664
x"fb0e0",-- -1266
x"f8dc0",-- -1828
x"f6aa0",-- -2390
x"f4bc0",-- -2884
x"f3470",-- -3257
x"f2640",-- -3484
x"f1d10",-- -3631
x"f1b10",-- -3663
x"f1fb0",-- -3589
x"f2c60",-- -3386
x"f4050",-- -3067
x"f5980",-- -2664
x"f7830",-- -2173
x"f9bf0",-- -1601
x"fc2a0",-- -982
x"fef00",-- -272
x"01680",-- 360
x"03e70",-- 999
x"06300",-- 1584
x"07b80",-- 1976
x"08ca0",-- 2250
x"09cc0",-- 2508
x"0a5e0",-- 2654
x"0a2a0",-- 2602
x"09e40",-- 2532
x"09880",-- 2440
x"08f20",-- 2290
x"07c40",-- 1988
x"06730",-- 1651
x"05240",-- 1316
x"03620",-- 866
x"01c60",-- 454
x"ffdb0",-- -37
x"fe340",-- -460
x"fcc10",-- -831
x"fb900",-- -1136
x"faca0",-- -1334
x"fa550",-- -1451
x"fa320",-- -1486
x"fa5d0",-- -1443
x"fad50",-- -1323
x"fb6c0",-- -1172
x"fc260",-- -986
x"fced0",-- -787
x"fd9c0",-- -612
x"fe3c0",-- -452
x"fef20",-- -270
x"ff710",-- -143
x"ffc20",-- -62
x"00120",-- 18
x"00940",-- 148
x"010b0",-- 267
x"01880",-- 392
x"02160",-- 534
x"02ef0",-- 751
x"03b70",-- 951
x"043c0",-- 1084
x"04e10",-- 1249
x"052b0",-- 1323
x"05540",-- 1364
x"054e0",-- 1358
x"05240",-- 1316
x"04db0",-- 1243
x"04a40",-- 1188
x"04a20",-- 1186
x"04fe0",-- 1278
x"05810",-- 1409
x"064e0",-- 1614
x"07a90",-- 1961
x"091f0",-- 2335
x"0acc0",-- 2764
x"0cf00",-- 3312
x"0f540",-- 3924
x"11720",-- 4466
x"12b90",-- 4793
x"13010",-- 4865
x"131d0",-- 4893
x"12370",-- 4663
x"10200",-- 4128
x"0ca20",-- 3234
x"091f0",-- 2335
x"06080",-- 1544
x"026e0",-- 622
x"fe570",-- -425
x"fabc0",-- -1348
x"f8960",-- -1898
x"f6480",-- -2488
x"f4250",-- -3035
x"f2350",-- -3531
x"f1200",-- -3808
x"f08c0",-- -3956
x"efbb0",-- -4165
x"ef8e0",-- -4210
x"ef880",-- -4216
x"efe70",-- -4121
x"f03c0",-- -4036
x"f1450",-- -3771
x"f2940",-- -3436
x"f3f30",-- -3085
x"f5a70",-- -2649
x"f7a20",-- -2142
x"fa200",-- -1504
x"fc710",-- -911
x"fe6c0",-- -404
x"003a0",-- 58
x"024d0",-- 589
x"03d00",-- 976
x"04a20",-- 1186
x"04dc0",-- 1244
x"04e10",-- 1249
x"049b0",-- 1179
x"03c40",-- 964
x"024b0",-- 587
x"00b20",-- 178
x"ff630",-- -157
x"fdc60",-- -570
x"fc340",-- -972
x"fad20",-- -1326
x"f98b0",-- -1653
x"f86c0",-- -1940
x"f7b70",-- -2121
x"f75e0",-- -2210
x"f7040",-- -2300
x"f7040",-- -2300
x"f74a0",-- -2230
x"f82a0",-- -2006
x"f9380",-- -1736
x"fa300",-- -1488
x"fb510",-- -1199
x"fcd40",-- -812
x"fe890",-- -375
x"ff6d0",-- -147
x"00280",-- 40
x"013f0",-- 319
x"02b70",-- 695
x"03cc0",-- 972
x"04340",-- 1076
x"05010",-- 1281
x"065f0",-- 1631
x"06f50",-- 1781
x"06980",-- 1688
x"06a40",-- 1700
x"066b0",-- 1643
x"05a40",-- 1444
x"04b80",-- 1208
x"03860",-- 902
x"029d0",-- 669
x"01d00",-- 464
x"00e40",-- 228
x"00620",-- 98
x"000a0",-- 10
x"ff7c0",-- -132
x"ff150",-- -235
x"ff580",-- -168
x"ff380",-- -200
x"ff220",-- -222
x"ff180",-- -232
x"fee60",-- -282
x"fefd0",-- -259
x"fef00",-- -272
x"fe370",-- -457
x"fe0c0",-- -500
x"fe550",-- -427
x"fe3f0",-- -449
x"fe5a0",-- -422
x"ff0e0",-- -242
x"ff8f0",-- -113
x"00110",-- 17
x"011c0",-- 284
x"013a0",-- 314
x"020f0",-- 527
x"02620",-- 610
x"02160",-- 534
x"02440",-- 580
x"02190",-- 537
x"02280",-- 552
x"01bd0",-- 445
x"02320",-- 562
x"02870",-- 647
x"02be0",-- 702
x"032c0",-- 812
x"039e0",-- 926
x"054f0",-- 1359
x"06690",-- 1641
x"07c90",-- 1993
x"094c0",-- 2380
x"0a930",-- 2707
x"0c280",-- 3112
x"0d710",-- 3441
x"0dbd0",-- 3517
x"0d360",-- 3382
x"0ce00",-- 3296
x"0c770",-- 3191
x"0b560",-- 2902
x"099e0",-- 2462
x"07bc0",-- 1980
x"06300",-- 1584
x"05010",-- 1281
x"02930",-- 659
x"008a0",-- 138
x"fec50",-- -315
x"fd5d0",-- -675
x"fc070",-- -1017
x"fa3f0",-- -1473
x"f8e80",-- -1816
x"f7810",-- -2175
x"f6580",-- -2472
x"f54f0",-- -2737
x"f4840",-- -2940
x"f3b30",-- -3149
x"f2c80",-- -3384
x"f3150",-- -3307
x"f3650",-- -3227
x"f3ea0",-- -3094
x"f4f80",-- -2824
x"f60c0",-- -2548
x"f7860",-- -2170
x"f9b20",-- -1614
x"fb600",-- -1184
x"fc4d0",-- -947
x"fe0a0",-- -502
x"ff710",-- -143
x"006b0",-- 107
x"01090",-- 265
x"01380",-- 312
x"011f0",-- 287
x"01220",-- 290
x"00f00",-- 240
x"00280",-- 40
x"ffb80",-- -72
x"ff110",-- -239
x"fe3e0",-- -450
x"fe0a0",-- -502
x"fd790",-- -647
x"fcd40",-- -812
x"fcbb0",-- -837
x"fcd50",-- -811
x"fcbb0",-- -837
x"fcf00",-- -784
x"fce60",-- -794
x"fd180",-- -744
x"fd7c0",-- -644
x"fe2d0",-- -467
x"fe660",-- -410
x"febb0",-- -325
x"ff860",-- -122
x"ffe90",-- -23
x"00bc0",-- 188
x"016f0",-- 367
x"01810",-- 385
x"01530",-- 339
x"018b0",-- 395
x"01940",-- 404
x"017e0",-- 382
x"01240",-- 292
x"007a0",-- 122
x"00c80",-- 200
x"01a60",-- 422
x"00f20",-- 242
x"00850",-- 133
x"01290",-- 297
x"014c0",-- 332
x"016a0",-- 362
x"01260",-- 294
x"01030",-- 259
x"012c0",-- 300
x"00c10",-- 193
x"01630",-- 355
x"010d0",-- 269
x"00cb0",-- 203
x"005a0",-- 90
x"00610",-- 97
x"00bc0",-- 188
x"ffdb0",-- -37
x"004b0",-- 75
x"ff8a0",-- -118
x"ffe70",-- -25
x"000a0",-- 10
x"fff60",-- -10
x"ffab0",-- -85
x"ffee0",-- -18
x"003a0",-- 58
x"ffcc0",-- -52
x"000c0",-- 12
x"fe3c0",-- -452
x"00bb0",-- 187
x"f8d50",-- -1835
x"fea20",-- -350
x"ff6c0",-- -148
x"f9130",-- -1773
x"01450",-- 325
x"fb310",-- -1231
x"ff420",-- -190
x"00250",-- 37
x"fd7c0",-- -644
x"013f0",-- 319
x"fe340",-- -460
x"00cb0",-- 203
x"01d50",-- 469
x"00000",-- 0
x"03c70",-- 967
x"03dd0",-- 989
x"044b0",-- 1099
x"05ec0",-- 1516
x"04990",-- 1177
x"06730",-- 1651
x"06480",-- 1608
x"072c0",-- 1836
x"07220",-- 1826
x"072c0",-- 1836
x"08bd0",-- 2237
x"08e50",-- 2277
x"094e0",-- 2382
x"09030",-- 2307
x"08ea0",-- 2282
x"07f40",-- 2036
x"07940",-- 1940
x"05d30",-- 1491
x"04bd0",-- 1213
x"04f20",-- 1266
x"03170",-- 791
x"01e40",-- 484
x"01590",-- 345
x"004b0",-- 75
x"ff8b0",-- -117
x"feaa0",-- -342
x"fe230",-- -477
x"fd680",-- -664
x"fbc40",-- -1084
x"fb450",-- -1211
x"fafd0",-- -1283
x"fa250",-- -1499
x"f90c0",-- -1780
x"f92c0",-- -1748
x"f9040",-- -1788
x"f8b40",-- -1868
x"f9700",-- -1680
x"f9c70",-- -1593
x"f9fd0",-- -1539
x"fad90",-- -1319
x"fc050",-- -1019
x"fc340",-- -972
x"fcac0",-- -852
x"fd760",-- -650
x"fd710",-- -655
x"fd970",-- -617
x"fd860",-- -634
x"fd530",-- -685
x"fcf70",-- -777
x"fd130",-- -749
x"fd4f0",-- -689
x"fcfc0",-- -772
x"fd560",-- -682
x"fd400",-- -704
x"fd530",-- -685
x"fdd50",-- -555
x"fe140",-- -492
x"fe260",-- -474
x"fe850",-- -379
x"ff060",-- -250
x"feff0",-- -257
x"ff5d0",-- -163
x"ffbd0",-- -67
x"ff510",-- -175
x"fff40",-- -12
x"ffe00",-- -32
x"00120",-- 18
x"00440",-- 68
x"fff10",-- -15
x"00de0",-- 222
x"008c0",-- 140
x"00f40",-- 244
x"00d90",-- 217
x"00e30",-- 227
x"01490",-- 329
x"017e0",-- 382
x"01a90",-- 425
x"01670",-- 359
x"01ea0",-- 490
x"01a90",-- 425
x"019a0",-- 410
x"01740",-- 372
x"012b0",-- 299
x"011f0",-- 287
x"00a80",-- 168
x"00d50",-- 213
x"00a50",-- 165
x"008e0",-- 142
x"007a0",-- 122
x"00bb0",-- 187
x"00da0",-- 218
x"00dc0",-- 220
x"00cf0",-- 207
x"00c00",-- 192
x"01060",-- 262
x"000f0",-- 15
x"00410",-- 65
x"001e0",-- 30
x"ffd60",-- -42
x"ff970",-- -105
x"feff0",-- -257
x"ff600",-- -160
x"fec80",-- -312
x"fed40",-- -300
x"fec10",-- -319
x"fe300",-- -464
x"fe730",-- -397
x"fe300",-- -464
x"fe2d0",-- -467
x"fe6e0",-- -402
x"fe3f0",-- -449
x"fe2a0",-- -470
x"fe430",-- -445
x"fe3c0",-- -452
x"feb90",-- -327
x"fed00",-- -304
x"ff4a0",-- -182
x"ff990",-- -103
x"ffad0",-- -83
x"00050",-- 5
x"fff80",-- -8
x"00760",-- 118
x"01180",-- 280
x"00e90",-- 233
x"00f40",-- 244
x"01f60",-- 502
x"01a90",-- 425
x"01ce0",-- 462
x"022f0",-- 559
x"025c0",-- 604
x"02940",-- 660
x"02710",-- 625
x"02fc0",-- 764
x"030e0",-- 782
x"033d0",-- 829
x"03650",-- 869
x"03c60",-- 966
x"04110",-- 1041
x"03da0",-- 986
x"04110",-- 1041
x"041b0",-- 1051
x"03e70",-- 999
x"03a10",-- 929
x"03b70",-- 951
x"036c0",-- 876
x"02f20",-- 754
x"02d60",-- 726
x"02a70",-- 679
x"026e0",-- 622
x"02250",-- 549
x"01ce0",-- 462
x"01b30",-- 435
x"01620",-- 354
x"00cf0",-- 207
x"007d0",-- 125
x"ffd60",-- -42
x"ff5b0",-- -165
x"fefc0",-- -260
x"fe350",-- -459
x"fdfe0",-- -514
x"fd7c0",-- -644
x"fd160",-- -746
x"fd310",-- -719
x"fcd00",-- -816
x"fcd00",-- -816
x"fcb10",-- -847
x"fcbb0",-- -837
x"fce10",-- -799
x"fce60",-- -794
x"fce30",-- -797
x"fca80",-- -856
x"fced0",-- -787
x"fcf00",-- -784
x"fcaa0",-- -854
x"fcaa0",-- -854
x"fc910",-- -879
x"fc780",-- -904
x"fc9e0",-- -866
x"fca50",-- -859
x"fc990",-- -871
x"fce30",-- -797
x"fceb0",-- -789
x"fd150",-- -747
x"fd530",-- -685
x"fd6c0",-- -660
x"fd8d0",-- -627
x"fdb80",-- -584
x"fde70",-- -537
x"fe1c0",-- -484
x"fe750",-- -395
x"fe9b0",-- -357
x"ff070",-- -249
x"ff800",-- -128
x"ffd10",-- -47
x"00260",-- 38
x"00870",-- 135
x"00d20",-- 210
x"01100",-- 272
x"01580",-- 344
x"01620",-- 354
x"01770",-- 375
x"01860",-- 390
x"018d0",-- 397
x"01a40",-- 420
x"01790",-- 377
x"01880",-- 392
x"01970",-- 407
x"01a40",-- 420
x"01a60",-- 422
x"018d0",-- 397
x"01a90",-- 425
x"018f0",-- 399
x"01860",-- 390
x"01830",-- 387
x"016a0",-- 362
x"01590",-- 345
x"01530",-- 339
x"01440",-- 324
x"01400",-- 320
x"01170",-- 279
x"00f50",-- 245
x"00eb0",-- 235
x"00b20",-- 178
x"00b90",-- 185
x"00800",-- 128
x"00640",-- 100
x"005d0",-- 93
x"00410",-- 65
x"003a0",-- 58
x"00210",-- 33
x"00160",-- 22
x"00120",-- 18
x"fffe0",-- -2
x"fffe0",-- -2
x"00050",-- 5
x"00000",-- 0
x"00020",-- 2
x"ffdf0",-- -33
x"fff40",-- -12
x"fff60",-- -10
x"fff90",-- -7
x"000d0",-- 13
x"00030",-- 3
x"00250",-- 37
x"00250",-- 37
x"00430",-- 67
x"004b0",-- 75
x"005d0",-- 93
x"00660",-- 102
x"00700",-- 112
x"008e0",-- 142
x"008f0",-- 143
x"00b90",-- 185
x"00c30",-- 195
x"00d50",-- 213
x"00eb0",-- 235
x"01090",-- 265
x"01260",-- 294
x"014e0",-- 334
x"01790",-- 377
x"01830",-- 387
x"01970",-- 407
x"01a90",-- 425
x"01a90",-- 425
x"01860",-- 390
x"01860",-- 390
x"015b0",-- 347
x"01380",-- 312
x"01290",-- 297
x"00dc0",-- 220
x"00a80",-- 168
x"00640",-- 100
x"002b0",-- 43
x"ffd80",-- -40
x"ff8d0",-- -115
x"ff290",-- -215
x"feeb0",-- -277
x"fea00",-- -352
x"fe490",-- -439
x"fe140",-- -492
x"fdc20",-- -574
x"fdab0",-- -597
x"fd6c0",-- -660
x"fd560",-- -682
x"fd4a0",-- -694
x"fd470",-- -697
x"fd530",-- -685
x"fd4a0",-- -694
x"fd560",-- -682
x"fd620",-- -670
x"fd710",-- -655
x"fd850",-- -635
x"fd920",-- -622
x"fdab0",-- -597
x"fdc10",-- -575
x"fdd00",-- -560
x"fe000",-- -512
x"fdf90",-- -519
x"fe070",-- -505
x"fe200",-- -480
x"fe1e0",-- -482
x"fe340",-- -460
x"fe430",-- -445
x"fe760",-- -394
x"fe890",-- -375
x"feaf0",-- -337
x"fee60",-- -282
x"ff240",-- -220
x"ff490",-- -183
x"ff6d0",-- -147
x"ffbd0",-- -67
x"fffe0",-- -2
x"00370",-- 55
x"004b0",-- 75
x"009d0",-- 157
x"00ed0",-- 237
x"01060",-- 262
x"013f0",-- 319
x"01310",-- 305
x"013b0",-- 315
x"01760",-- 374
x"01710",-- 369
x"01900",-- 400
x"01b50",-- 437
x"01e20",-- 482
x"01c10",-- 449
x"01db0",-- 475
x"02000",-- 512
x"01f40",-- 500
x"02030",-- 515
x"01c70",-- 455
x"01db0",-- 475
x"01c70",-- 455
x"01cc0",-- 460
x"019e0",-- 414
x"01710",-- 369
x"01680",-- 360
x"01490",-- 329
x"01100",-- 272
x"00d40",-- 212
x"00b90",-- 185
x"00800",-- 128
x"00990",-- 153
x"006c0",-- 108
x"003f0",-- 63
x"00320",-- 50
x"00200",-- 32
x"00080",-- 8
x"fff40",-- -12
x"ffdf0",-- -33
x"ffc60",-- -58
x"ffc60",-- -58
x"ffa90",-- -87
x"ff990",-- -103
x"ff710",-- -143
x"ff650",-- -155
x"ff4a0",-- -182
x"ff4e0",-- -178
x"ff3b0",-- -197
x"ff350",-- -203
x"ff1f0",-- -225
x"ff170",-- -233
x"ff270",-- -217
x"ff260",-- -218
x"ff1f0",-- -225
x"ff180",-- -232
x"ff2e0",-- -210
x"ff290",-- -215
x"ff560",-- -170
x"ff580",-- -168
x"ff850",-- -123
x"ff8a0",-- -118
x"ff900",-- -112
x"ffbc0",-- -68
x"ffcc0",-- -52
x"fff30",-- -13
x"000d0",-- 13
x"00260",-- 38
x"00410",-- 65
x"006b0",-- 107
x"00930",-- 147
x"00b90",-- 185
x"00e10",-- 225
x"00f90",-- 249
x"010d0",-- 269
x"012e0",-- 302
x"01310",-- 305
x"01310",-- 305
x"012c0",-- 300
x"012e0",-- 302
x"01300",-- 304
x"012e0",-- 302
x"01180",-- 280
x"00fc0",-- 252
x"01010",-- 257
x"00ed0",-- 237
x"00e60",-- 230
x"00e40",-- 228
x"00d20",-- 210
x"00de0",-- 222
x"00cb0",-- 203
x"00ac0",-- 172
x"009d0",-- 157
x"00750",-- 117
x"005d0",-- 93
x"00440",-- 68
x"002b0",-- 43
x"00000",-- 0
x"ffd10",-- -47
x"ffb80",-- -72
x"ff8b0",-- -117
x"ff710",-- -143
x"ff4a0",-- -182
x"ff330",-- -205
x"ff150",-- -235
x"ff070",-- -249
x"feee0",-- -274
x"feed0",-- -275
x"feda0",-- -294
x"fec50",-- -315
x"fedc0",-- -292
x"feaf0",-- -337
x"fec10",-- -319
x"feb20",-- -334
x"feac0",-- -340
x"feb60",-- -330
x"fead0",-- -339
x"feca0",-- -310
x"feca0",-- -310
x"fef50",-- -267
x"fefd0",-- -259
x"ff210",-- -223
x"ff420",-- -190
x"ff560",-- -170
x"ff600",-- -160
x"ff850",-- -123
x"ff720",-- -142
x"ff8a0",-- -118
x"001b0",-- 27
x"ffda0",-- -38
x"ffea0",-- -22
x"fff10",-- -15
x"00030",-- 3
x"00460",-- 70
x"00480",-- 72
x"00750",-- 117
x"00730",-- 115
x"00910",-- 145
x"00a00",-- 160
x"00cb0",-- 203
x"00250",-- 37
x"fe8a0",-- -374
x"fdee0",-- -530
x"feee0",-- -274
x"000c0",-- 12
x"00e80",-- 232
x"01450",-- 325
x"00f90",-- 249
x"01310",-- 305
x"01130",-- 275
x"00c10",-- 193
x"00ac0",-- 172
x"00730",-- 115
x"008e0",-- 142
x"00c80",-- 200
x"012b0",-- 299
x"015b0",-- 347
x"01c90",-- 457
x"01e70",-- 487
x"01b50",-- 437
x"01650",-- 357
x"00f90",-- 249
x"00df0",-- 223
x"00be0",-- 190
x"00df0",-- 223
x"007b0",-- 123
x"00410",-- 65
x"00120",-- 18
x"ffce0",-- -50
x"00460",-- 70
x"005a0",-- 90
x"000c0",-- 12
x"fff90",-- -7
x"001e0",-- 30
x"004b0",-- 75
x"002d0",-- 45
x"002f0",-- 47
x"00000",-- 0
x"00080",-- 8
x"fff60",-- -10
x"fff40",-- -12
x"ffe90",-- -23
x"ffdf0",-- -33
x"ffe70",-- -25
x"ffdb0",-- -37
x"ffe50",-- -27
x"ff9c0",-- -100
x"ffab0",-- -85
x"ffa60",-- -90
x"ffa80",-- -88
x"ffcc0",-- -52
x"ff950",-- -107
x"ff830",-- -125
x"ff7e0",-- -130
x"ff790",-- -135
x"ff920",-- -110
x"ff8b0",-- -117
x"ff8a0",-- -118
x"ff800",-- -128
x"ff8d0",-- -115
x"ffa90",-- -87
x"ff900",-- -112
x"ff810",-- -127
x"ff6f0",-- -145
x"ff790",-- -135
x"ff830",-- -125
x"ff9c0",-- -100
x"ff760",-- -138
x"ff670",-- -153
x"ff7e0",-- -130
x"ff5d0",-- -163
x"ff720",-- -142
x"ff600",-- -160
x"ff330",-- -205
x"ff680",-- -152
x"ff630",-- -157
x"ff560",-- -170
x"ff590",-- -167
x"ff470",-- -185
x"ff530",-- -173
x"ff380",-- -200
x"ff8a0",-- -118
x"ff350",-- -203
x"ff710",-- -143
x"ff630",-- -157
x"ff420",-- -190
x"ff9c0",-- -100
x"ff1c0",-- -228
x"ff5d0",-- -163
x"ff6a0",-- -150
x"ff670",-- -153
x"ff830",-- -125
x"ff770",-- -137
x"ff5d0",-- -163
x"ff810",-- -127
x"ff6d0",-- -147
x"ff6f0",-- -145
x"ffad0",-- -83
x"ff860",-- -122
x"ffce0",-- -50
x"ffa30",-- -93
x"ffe50",-- -27
x"fff80",-- -8
x"00170",-- 23
x"00000",-- 0
x"00070",-- 7
x"00410",-- 65
x"002a0",-- 42
x"006b0",-- 107
x"001e0",-- 30
x"00520",-- 82
x"004b0",-- 75
x"005d0",-- 93
x"00a00",-- 160
x"00640",-- 100
x"00980",-- 152
x"00800",-- 128
x"00870",-- 135
x"00a30",-- 163
x"00ac0",-- 172
x"00890",-- 137
x"00d70",-- 215
x"00bc0",-- 188
x"00e80",-- 232
x"00df0",-- 223
x"00930",-- 147
x"01010",-- 257
x"00960",-- 150
x"00eb0",-- 235
x"00e60",-- 230
x"00d70",-- 215
x"00dc0",-- 220
x"011f0",-- 287
x"00cb0",-- 203
x"013b0",-- 315
x"00d50",-- 213
x"011c0",-- 284
x"01450",-- 325
x"00af0",-- 175
x"01240",-- 292
x"00a30",-- 163
x"00d50",-- 213
x"00af0",-- 175
x"009d0",-- 157
x"008f0",-- 143
x"006b0",-- 107
x"00710",-- 113
x"00490",-- 73
x"007b0",-- 123
x"00620",-- 98
x"00430",-- 67
x"00640",-- 100
x"00350",-- 53
x"00000",-- 0
x"00410",-- 65
x"ffe50",-- -27
x"ffcc0",-- -52
x"ffee0",-- -18
x"ffa90",-- -87
x"fffb0",-- -5
x"000f0",-- 15
x"00070",-- 7
x"fff40",-- -12
x"00050",-- 5
x"ffda0",-- -38
x"fffb0",-- -5
x"ffdf0",-- -33
x"ffd80",-- -40
x"ffc60",-- -58
x"ffc90",-- -55
x"ffb50",-- -75
x"ff8a0",-- -118
x"ffb70",-- -73
x"ff710",-- -143
x"ff600",-- -160
x"ff800",-- -128
x"ff800",-- -128
x"ff800",-- -128
x"ffad0",-- -83
x"ff900",-- -112
x"ff830",-- -125
x"ff580",-- -168
x"ff6a0",-- -150
x"ff6d0",-- -147
x"ff7c0",-- -132
x"ff830",-- -125
x"ff560",-- -170
x"ff630",-- -157
x"ff4a0",-- -182
x"ff790",-- -135
x"ff510",-- -175
x"ff5e0",-- -162
x"ff5d0",-- -163
x"ff600",-- -160
x"ff2c0",-- -212
x"ff2e0",-- -210
x"ff6a0",-- -150
x"ff470",-- -185
x"ff400",-- -192
x"ff7b0",-- -133
x"ff810",-- -127
x"ff540",-- -172
x"ff900",-- -112
x"ff6c0",-- -148
x"ff6d0",-- -147
x"ff950",-- -107
x"ff310",-- -207
x"ff7b0",-- -133
x"ff600",-- -160
x"ff3d0",-- -195
x"ff970",-- -105
x"ff950",-- -107
x"ffae0",-- -82
x"ffe70",-- -25
x"ffa60",-- -90
x"ffae0",-- -82
x"ffc20",-- -62
x"ff800",-- -128
x"ff950",-- -107
x"ff970",-- -105
x"ffbc0",-- -68
x"ffe40",-- -28
x"ffa60",-- -90
x"ffec0",-- -20
x"ffea0",-- -22
x"ffe20",-- -30
x"00120",-- 18
x"00170",-- 23
x"00210",-- 33
x"fff40",-- -12
x"005a0",-- 90
x"ffe20",-- -30
x"00530",-- 83
x"006c0",-- 108
x"00200",-- 32
x"00370",-- 55
x"00000",-- 0
x"00930",-- 147
x"00210",-- 33
x"00700",-- 112
x"00640",-- 100
x"00250",-- 37
x"00370",-- 55
x"fffd0",-- -3
x"00670",-- 103
x"00da0",-- 218
x"00c30",-- 195
x"00fc0",-- 252
x"00f90",-- 249
x"00e80",-- 232
x"00b90",-- 185
x"00840",-- 132
x"00610",-- 97
x"00930",-- 147
x"00ad0",-- 173
x"003a0",-- 58
x"003e0",-- 62
x"00120",-- 18
x"002a0",-- 42
x"00850",-- 133
x"004b0",-- 75
x"007a0",-- 122
x"00480",-- 72
x"00c10",-- 193
x"00760",-- 118
x"00730",-- 115
x"00000",-- 0
x"000f0",-- 15
x"00110",-- 17
x"ffea0",-- -22
x"005f0",-- 95
x"ffb20",-- -78
x"00640",-- 100
x"00960",-- 150
x"00a50",-- 165
x"00390",-- 57
x"fff90",-- -7
x"00120",-- 18
x"00370",-- 55
x"00840",-- 132
x"ffc20",-- -62
x"ff4e0",-- -178
x"00080",-- 8
x"00080",-- 8
x"ffa40",-- -92
x"000c0",-- 12
x"ffe50",-- -27
x"ff740",-- -140
x"ff710",-- -143
x"ff900",-- -112
x"00160",-- 22
x"ff830",-- -125
x"ffc70",-- -57
x"ffe40",-- -28
x"ffb30",-- -77
x"ffa60",-- -90
x"ffb50",-- -75
x"ff650",-- -155
x"ff5b0",-- -165
x"ffe00",-- -32
x"fee60",-- -282
x"ff450",-- -187
x"ffd60",-- -42
x"ffd10",-- -47
x"ffbf0",-- -65
x"ff850",-- -123
x"fee80",-- -280
x"ff2c0",-- -212
x"ff990",-- -103
x"ff350",-- -203
x"fee10",-- -287
x"ff4c0",-- -180
x"ffe20",-- -30
x"ff630",-- -157
x"ffef0",-- -17
x"fff10",-- -15
x"ff630",-- -157
x"00020",-- 2
x"ff670",-- -153
x"ff1f0",-- -225
x"ffc20",-- -62
x"00320",-- 50
x"ffc20",-- -62
x"ffa40",-- -92
x"004e0",-- 78
x"ff8d0",-- -115
x"ffa10",-- -95
x"ff900",-- -112
x"ff490",-- -183
x"001e0",-- 30
x"ffdf0",-- -33
x"ffe50",-- -27
x"ff4a0",-- -182
x"ffec0",-- -20
x"00430",-- 67
x"ff580",-- -168
x"00200",-- 32
x"ffe20",-- -30
x"ffe20",-- -30
x"ffc60",-- -58
x"ffa30",-- -93
x"00c30",-- 195
x"ffd50",-- -43
x"006b0",-- 107
x"00d40",-- 212
x"00250",-- 37
x"00610",-- 97
x"00700",-- 112
x"00c30",-- 195
x"004e0",-- 78
x"00960",-- 150
x"00250",-- 37
x"00500",-- 80
x"ffad0",-- -83
x"00530",-- 83
x"007d0",-- 125
x"00fe0",-- 254
x"01260",-- 294
x"ff540",-- -172
x"ffdd0",-- -35
x"002a0",-- 42
x"01180",-- 280
x"01860",-- 390
x"00ac0",-- 172
x"01c20",-- 450
x"01770",-- 375
x"007b0",-- 123
x"fff40",-- -12
x"00700",-- 112
x"01ad0",-- 429
x"00120",-- 18
x"007f0",-- 127
x"00e60",-- 230
x"00120",-- 18
x"008a0",-- 138
x"006c0",-- 108
x"003e0",-- 62
x"ffee0",-- -18
x"00570",-- 87
x"000f0",-- 15
x"00200",-- 32
x"ffc90",-- -55
x"001b0",-- 27
x"00210",-- 33
x"002a0",-- 42
x"005a0",-- 90
x"00440",-- 68
x"01210",-- 289
x"01600",-- 352
x"01710",-- 369
x"00e80",-- 232
x"005a0",-- 90
x"ff540",-- -172
x"feed0",-- -275
x"ff590",-- -167
x"ffc60",-- -58
x"ffb20",-- -78
x"ffdf0",-- -33
x"00800",-- 128
x"00f50",-- 245
x"ffd30",-- -45
x"ff270",-- -217
x"fe520",-- -430
x"fe0d0",-- -499
x"ff040",-- -252
x"feaa0",-- -342
x"ff710",-- -143
x"ffa80",-- -88
x"009d0",-- 157
x"00ff0",-- 255
x"ffbc0",-- -68
x"fee60",-- -282
x"fdce0",-- -562
x"fdda0",-- -550
x"fe570",-- -425
x"fde90",-- -535
x"ff180",-- -232
x"00550",-- 85
x"00ca0",-- 202
x"002b0",-- 43
x"fff80",-- -8
x"ff490",-- -183
x"fdfe0",-- -514
x"fdb80",-- -584
x"fd740",-- -652
x"fe350",-- -459
x"fe160",-- -490
x"ff150",-- -235
x"ffbf0",-- -65
x"ffa10",-- -95
x"ffd30",-- -45
x"ffa80",-- -88
x"ff5e0",-- -162
x"fe960",-- -362
x"fea80",-- -344
x"ff010",-- -255
x"ff270",-- -217
x"ff0e0",-- -242
x"00440",-- 68
x"00be0",-- 190
x"00ff0",-- 255
x"fec80",-- -312
x"fd330",-- -717
x"fb740",-- -1164
x"f8f20",-- -1806
x"fa550",-- -1451
x"fbf30",-- -1037
x"fe4b0",-- -437
x"00390",-- 57
x"01bf0",-- 447
x"03830",-- 899
x"03ee0",-- 1006
x"03940",-- 916
x"02e80",-- 744
x"02430",-- 579
x"024b0",-- 587
x"01850",-- 389
x"03360",-- 822
x"03300",-- 816
x"04660",-- 1126
x"05760",-- 1398
x"05470",-- 1351
x"05770",-- 1399
x"043a0",-- 1082
x"03880",-- 904
x"02320",-- 562
x"01d50",-- 469
x"00520",-- 82
x"ff3a0",-- -198
x"fef80",-- -264
x"ff3a0",-- -198
x"ffae0",-- -82
x"ff830",-- -125
x"00000",-- 0
x"ff740",-- -140
x"ffdf0",-- -33
x"013f0",-- 319
x"01060",-- 262
x"00dc0",-- 220
x"008f0",-- 143
x"01510",-- 337
x"01810",-- 385
x"01b30",-- 435
x"018f0",-- 399
x"01060",-- 262
x"025f0",-- 607
x"02000",-- 512
x"01450",-- 325
x"00890",-- 137
x"00280",-- 40
x"00ad0",-- 173
x"00f20",-- 242
x"00f90",-- 249
x"00a80",-- 168
x"00f90",-- 249
x"01e00",-- 480
x"026b0",-- 619
x"01dd0",-- 477
x"000c0",-- 12
x"ffa30",-- -93
x"fe490",-- -439
x"fe1e0",-- -482
x"fe3f0",-- -449
x"fd530",-- -685
x"fd0c0",-- -756
x"fdda0",-- -550
x"fe1b0",-- -485
x"fe570",-- -425
x"fe170",-- -489
x"f98b0",-- -1653
x"fe890",-- -375
x"fbc90",-- -1079
x"fd3a0",-- -710
x"fff30",-- -13
x"fc1c0",-- -996
x"00210",-- 33
x"febb0",-- -325
x"fe5c0",-- -420
x"fe5d0",-- -419
x"fd800",-- -640
x"fe140",-- -492
x"fe570",-- -425
x"ff790",-- -135
x"ffc70",-- -57
x"fee40",-- -284
x"ff8b0",-- -117
x"feda0",-- -294
x"fedf0",-- -289
x"ff0e0",-- -242
x"fd4e0",-- -690
x"fdf80",-- -520
x"fce60",-- -794
x"fcfc0",-- -772
x"fd3b0",-- -709
x"fd2e0",-- -722
x"fd0c0",-- -756
x"fd760",-- -650
x"fe5a0",-- -422
x"fe190",-- -487
x"ff400",-- -192
x"ff0e0",-- -242
x"ff0c0",-- -244
x"ffbf0",-- -65
x"ff3b0",-- -197
x"ff6a0",-- -150
x"00070",-- 7
x"ffb00",-- -80
x"00ed0",-- 237
x"007f0",-- 127
x"011a0",-- 282
x"012b0",-- 299
x"016a0",-- 362
x"02020",-- 514
x"01030",-- 259
x"00f00",-- 240
x"00a00",-- 160
x"01600",-- 352
x"01450",-- 325
x"01620",-- 354
x"028a0",-- 650
x"01c10",-- 449
x"02550",-- 597
x"033b0",-- 827
x"03b00",-- 944
x"04710",-- 1137
x"04170",-- 1047
x"04080",-- 1032
x"04a20",-- 1186
x"05a40",-- 1444
x"073f0",-- 1855
x"08160",-- 2070
x"08e00",-- 2272
x"0a520",-- 2642
x"0ae80",-- 2792
x"0c2d0",-- 3117
x"0cd20",-- 3282
x"0d080",-- 3336
x"0df30",-- 3571
x"0e700",-- 3696
x"0fce0",-- 4046
x"0f920",-- 3986
x"0e540",-- 3668
x"0cae0",-- 3246
x"096a0",-- 2410
x"07800",-- 1920
x"04110",-- 1041
x"007a0",-- 122
x"fdd30",-- -557
x"fb6d0",-- -1171
x"fb110",-- -1263
x"f9570",-- -1705
x"f7ce0",-- -2098
x"f5ba0",-- -2630
x"f32c0",-- -3284
x"f1590",-- -3751
x"eeb40",-- -4428
x"ecfc0",-- -4868
x"eadf0",-- -5409
x"ea880",-- -5496
x"ec370",-- -5065
x"eeb90",-- -4423
x"f1d80",-- -3624
x"f4280",-- -3032
x"f74f0",-- -2225
x"fa640",-- -1436
x"fd650",-- -667
x"ff950",-- -107
x"007a0",-- 122
x"01c90",-- 457
x"032c0",-- 812
x"04b80",-- 1208
x"06020",-- 1538
x"06b10",-- 1713
x"06d20",-- 1746
x"06cd0",-- 1741
x"06c30",-- 1731
x"059a0",-- 1434
x"039a0",-- 922
x"01060",-- 262
x"febe0",-- -322
x"fced0",-- -787
x"fb430",-- -1213
x"f96b0",-- -1685
x"f7880",-- -2168
x"f6660",-- -2458
x"f4120",-- -3054
x"f30e0",-- -3314
x"f14a0",-- -3766
x"ef860",-- -4218
x"ed970",-- -4713
x"ed290",-- -4823
x"ee490",-- -4535
x"efef0",-- -4113
x"f1790",-- -3719
x"f3b00",-- -3152
x"f7920",-- -2158
x"fa6c0",-- -1428
x"fce10",-- -799
x"fe5f0",-- -417
x"ffdb0",-- -37
x"00cd0",-- 205
x"02910",-- 657
x"04760",-- 1142
x"06390",-- 1593
x"077b0",-- 1915
x"091f0",-- 2335
x"0a7a0",-- 2682
x"0b630",-- 2915
x"0a8e0",-- 2702
x"08f70",-- 2295
x"072c0",-- 1836
x"05560",-- 1366
x"03c40",-- 964
x"02370",-- 567
x"01580",-- 344
x"00580",-- 88
x"ffc60",-- -58
x"ffee0",-- -18
x"ff990",-- -103
x"febe0",-- -322
x"fdea0",-- -534
x"fdb30",-- -589
x"ff010",-- -255
x"ffcc0",-- -52
x"016d0",-- 365
x"03fe0",-- 1022
x"07350",-- 1845
x"0a190",-- 2585
x"0d290",-- 3369
x"0f760",-- 3958
x"127c0",-- 4732
x"144a0",-- 5194
x"15ce0",-- 5582
x"18540",-- 6228
x"1a2a0",-- 6698
x"1c9a0",-- 7322
x"1cd30",-- 7379
x"1d640",-- 7524
x"1ee50",-- 7909
x"1d5d0",-- 7517
x"19420",-- 6466
x"12400",-- 4672
x"0dc40",-- 3524
x"073f0",-- 1855
x"00a50",-- 165
x"fc020",-- -1022
x"f7c70",-- -2105
x"f5610",-- -2719
x"f1860",-- -3706
x"efde0",-- -4130
x"ed8e0",-- -4722
x"e9570",-- -5801
x"e4030",-- -7165
x"e0940",-- -8044
x"df730",-- -8333
x"de300",-- -8656
x"df540",-- -8364
x"e3650",-- -7323
x"e8c10",-- -5951
x"ef720",-- -4238
x"f59a0",-- -2662
x"fb330",-- -1229
x"ff9f0",-- -97
x"03300",-- 816
x"05e90",-- 1513
x"08ac0",-- 2220
x"0bf90",-- 3065
x"0dcb0",-- 3531
x"0ffa0",-- 4090
x"13580",-- 4952
x"15450",-- 5445
x"14980",-- 5272
x"12870",-- 4743
x"0f830",-- 3971
x"0b590",-- 2905
x"06a90",-- 1705
x"017e0",-- 382
x"fd6d0",-- -659
x"f9ec0",-- -1556
x"f67b0",-- -2437
x"f4580",-- -2984
x"f2870",-- -3449
x"efc40",-- -4156
x"ec300",-- -5072
x"e9970",-- -5737
x"e8000",-- -6144
x"e6990",-- -6503
x"e6530",-- -6573
x"e7d60",-- -6186
x"eac00",-- -5440
x"ef740",-- -4236
x"f3b60",-- -3146
x"f83a0",-- -1990
x"fbf90",-- -1031
x"fe390",-- -455
x"ffad0",-- -83
x"01e00",-- 480
x"04af0",-- 1199
x"05c70",-- 1479
x"07540",-- 1876
x"09040",-- 2308
x"0b350",-- 2869
x"0c410",-- 3137
x"0cb60",-- 3254
x"0c500",-- 3152
x"0a720",-- 2674
x"07bf0",-- 1983
x"051f0",-- 1311
x"03b80",-- 952
x"013b0",-- 315
x"feff0",-- -257
x"fd1a0",-- -742
x"fc230",-- -989
x"fb620",-- -1182
x"f9830",-- -1661
x"f8580",-- -1960
x"f7470",-- -2233
x"f66c0",-- -2452
x"f6a50",-- -2395
x"f7290",-- -2263
x"f8800",-- -1920
x"fa760",-- -1418
x"fc050",-- -1019
x"fe5c0",-- -420
x"00eb0",-- 235
x"02260",-- 550
x"02fe0",-- 766
x"046c0",-- 1132
x"05c20",-- 1474
x"072b0",-- 1835
x"085e0",-- 2142
x"0a230",-- 2595
x"0c690",-- 3177
x"0d900",-- 3472
x"0f3b0",-- 3899
x"103c0",-- 4156
x"10a20",-- 4258
x"10b90",-- 4281
x"10db0",-- 4315
x"12090",-- 4617
x"11b90",-- 4537
x"115d0",-- 4445
x"12bb0",-- 4795
x"14ca0",-- 5322
x"16db0",-- 5851
x"17f80",-- 6136
x"17d50",-- 6101
x"17e40",-- 6116
x"173f0",-- 5951
x"13b20",-- 5042
x"0c220",-- 3106
x"05b00",-- 1456
x"fef00",-- -272
x"f9ef0",-- -1553
x"f8000",-- -2048
x"f5250",-- -2779
x"f4850",-- -2939
x"f1d40",-- -3628
x"efec0",-- -4116
x"ee910",-- -4463
x"ea6e0",-- -5522
x"e3f40",-- -7180
x"df720",-- -8334
x"dfc50",-- -8251
x"e11b0",-- -7909
x"e39f0",-- -7265
x"e9d80",-- -5672
x"efbf0",-- -4161
x"f4e90",-- -2839
x"fa5c0",-- -1444
x"fe5a0",-- -422
x"00570",-- 87
x"020a0",-- 522
x"04d40",-- 1236
x"08c20",-- 2242
x"0e4b0",-- 3659
x"11f10",-- 4593
x"135d0",-- 4957
x"151d0",-- 5405
x"14bd0",-- 5309
x"11440",-- 4420
x"0bfe0",-- 3070
x"06280",-- 1576
x"00be0",-- 190
x"fd160",-- -746
x"fab10",-- -1359
x"f8ee0",-- -1810
x"f7450",-- -2235
x"f4140",-- -3052
x"f1200",-- -3808
x"ee820",-- -4478
x"ea8d0",-- -5491
x"e6100",-- -6640
x"e39d0",-- -7267
x"e3bf0",-- -7233
x"e5790",-- -6791
x"e8880",-- -6008
x"ecd50",-- -4907
x"efe30",-- -4125
x"f3310",-- -3279
x"f5da0",-- -2598
x"f8d40",-- -1836
x"fbbd0",-- -1091
x"fe350",-- -459
x"02210",-- 545
x"05b20",-- 1458
x"0bda0",-- 3034
x"0ee30",-- 3811
x"10250",-- 4133
x"11450",-- 4421
x"0feb0",-- 4075
x"0f1a0",-- 3866
x"0cf90",-- 3321
x"0b150",-- 2837
x"09c70",-- 2503
x"08580",-- 2136
x"07ce0",-- 1998
x"065d0",-- 1629
x"040a0",-- 1034
x"00e60",-- 230
x"fd3a0",-- -710
x"fa1e0",-- -1506
x"f7ab0",-- -2133
x"f5930",-- -2669
x"f4e90",-- -2839
x"f51a0",-- -2790
x"f5bd0",-- -2627
x"f7220",-- -2270
x"f84e0",-- -1970
x"f8410",-- -1983
x"f93e0",-- -1730
x"fa1e0",-- -1506
x"fc4d0",-- -947
x"fe620",-- -414
x"00840",-- 132
x"03360",-- 822
x"05360",-- 1334
x"07e40",-- 2020
x"082f0",-- 2095
x"09580",-- 2392
x"09c60",-- 2502
x"0a860",-- 2694
x"0cac0",-- 3244
x"0e4a0",-- 3658
x"100f0",-- 4111
x"10b30",-- 4275
x"118d0",-- 4493
x"120f0",-- 4623
x"12c00",-- 4800
x"11900",-- 4496
x"104f0",-- 4175
x"11800",-- 4480
x"12220",-- 4642
x"151c0",-- 5404
x"162f0",-- 5679
x"18140",-- 6164
x"18f90",-- 6393
x"17970",-- 6039
x"187a0",-- 6266
x"11090",-- 4361
x"07030",-- 1795
x"014e0",-- 334
x"faa00",-- -1376
x"f86b0",-- -1941
x"f57e0",-- -2690
x"f20b0",-- -3573
x"f0a20",-- -3934
x"ee7d0",-- -4483
x"eded0",-- -4627
x"ec760",-- -5002
x"e7ca0",-- -6198
x"dfe20",-- -8222
x"dd430",-- -8893
x"e0560",-- -8106
x"e4010",-- -7167
x"e8510",-- -6063
x"ee190",-- -4583
x"f3420",-- -3262
x"f84b0",-- -1973
x"fe5d0",-- -419
x"005d0",-- 93
x"01290",-- 297
x"049b0",-- 1179
x"08280",-- 2088
x"0e1d0",-- 3613
x"14820",-- 5250
x"16160",-- 5654
x"15820",-- 5506
x"15440",-- 5444
x"129d0",-- 4765
x"0d310",-- 3377
x"06930",-- 1683
x"00730",-- 115
x"fccf0",-- -817
x"fba60",-- -1114
x"fa350",-- -1483
x"f83f0",-- -1985
x"f48e0",-- -2930
x"efce0",-- -4146
x"ec370",-- -5065
x"e9a90",-- -5719
x"e5e50",-- -6683
x"e2f30",-- -7437
x"e35e0",-- -7330
x"e7180",-- -6376
x"eb040",-- -5372
x"ef2e0",-- -4306
x"f1970",-- -3689
x"f3ba0",-- -3142
x"f4f70",-- -2825
x"f4780",-- -2952
x"f95c0",-- -1700
x"fdec0",-- -532
x"03fd0",-- 1021
x"080c0",-- 2060
x"0ce10",-- 3297
x"14140",-- 5140
x"14250",-- 5157
x"11090",-- 4361
x"0ffd0",-- 4093
x"0e4d0",-- 3661
x"0c310",-- 3121
x"0bd80",-- 3032
x"0b120",-- 2834
x"0b400",-- 2880
x"09ad0",-- 2477
x"07090",-- 1801
x"047f0",-- 1151
x"fee90",-- -279
x"f97e0",-- -1666
x"f5f30",-- -2573
x"f5160",-- -2794
x"f6140",-- -2540
x"f6250",-- -2523
x"f6390",-- -2503
x"f78e0",-- -2162
x"f6f70",-- -2313
x"f60c0",-- -2548
x"f6000",-- -2560
x"f5920",-- -2670
x"f8250",-- -2011
x"fad50",-- -1323
x"fef80",-- -264
x"04a50",-- 1189
x"067f0",-- 1663
x"07220",-- 1826
x"07e90",-- 2025
x"08840",-- 2180
x"07cb0",-- 1995
x"080c0",-- 2060
x"09f90",-- 2553
x"0cc70",-- 3271
x"0f510",-- 3921
x"11680",-- 4456
x"12b80",-- 4792
x"11a60",-- 4518
x"10590",-- 4185
x"0ed20",-- 3794
x"0fc10",-- 4033
x"10fa0",-- 4346
x"0f620",-- 3938
x"11680",-- 4456
x"13150",-- 4885
x"166d0",-- 5741
x"17420",-- 5954
x"15dd0",-- 5597
x"15e90",-- 5609
x"13f80",-- 5112
x"14630",-- 5219
x"0d5b0",-- 3419
x"05a40",-- 1444
x"fd710",-- -655
x"f60f0",-- -2545
x"f6ca0",-- -2358
x"f6120",-- -2542
x"f4550",-- -2987
x"ef7f0",-- -4225
x"ec640",-- -5020
x"eb560",-- -5290
x"e96d0",-- -5779
x"e4100",-- -7152
x"ddc90",-- -8759
x"ddf70",-- -8713
x"e1f10",-- -7695
x"e7660",-- -6298
x"edba0",-- -4678
x"f2910",-- -3439
x"f3f80",-- -3080
x"f7380",-- -2248
x"fce60",-- -794
x"ff8d0",-- -115
x"01e00",-- 480
x"05fe0",-- 1534
x"0bd80",-- 3032
x"139b0",-- 5019
x"18cc0",-- 6348
x"17b00",-- 6064
x"146b0",-- 5227
x"119a0",-- 4506
x"0d3d0",-- 3389
x"09740",-- 2420
x"06700",-- 1648
x"01f90",-- 505
x"ff060",-- -250
x"fe6b0",-- -405
x"fc910",-- -879
x"f7b80",-- -2120
x"f0e10",-- -3871
x"e9c40",-- -5692
x"e6dd0",-- -6435
x"e6b20",-- -6478
x"e6380",-- -6600
x"e6330",-- -6605
x"e7fb0",-- -6149
x"ea140",-- -5612
x"ebf70",-- -5129
x"eecb0",-- -4405
x"ef100",-- -4336
x"ef2e0",-- -4306
x"efa60",-- -4186
x"f4c60",-- -2874
x"fdec0",-- -532
x"05470",-- 1351
x"09f10",-- 2545
x"0bb30",-- 2995
x"0fbd0",-- 4029
x"120e0",-- 4622
x"104b0",-- 4171
x"0f220",-- 3874
x"0f060",-- 3846
x"0f380",-- 3896
x"10cd0",-- 4301
x"12720",-- 4722
x"10af0",-- 4271
x"0c220",-- 3106
x"06a20",-- 1698
x"02c60",-- 710
x"ff6d0",-- -147
x"fb510",-- -1199
x"f8cf0",-- -1841
x"f7a40",-- -2140
x"f8c00",-- -1856
x"f9340",-- -1740
x"f6b10",-- -2383
x"f43c0",-- -3012
x"f15b0",-- -3749
x"efde0",-- -4130
x"f2120",-- -3566
x"f5150",-- -2795
x"f86c0",-- -1940
x"fb200",-- -1248
x"fe500",-- -432
x"02610",-- 609
x"04260",-- 1062
x"03530",-- 851
x"036c0",-- 876
x"05df0",-- 1503
x"09290",-- 2345
x"0c6e0",-- 3182
x"0efe0",-- 3838
x"10d60",-- 4310
x"10660",-- 4198
x"10610",-- 4193
x"10b30",-- 4275
x"0f180",-- 3864
x"0e040",-- 3588
x"0d990",-- 3481
x"0f3d0",-- 3901
x"12f20",-- 4850
x"12540",-- 4692
x"11680",-- 4456
x"0f560",-- 3926
x"0e930",-- 3731
x"10250",-- 4133
x"0fab0",-- 4011
x"12930",-- 4755
x"12900",-- 4752
x"13a10",-- 5025
x"15360",-- 5430
x"0f940",-- 3988
x"06b40",-- 1716
x"fadf0",-- -1313
x"f4a00",-- -2912
x"f62a0",-- -2518
x"f7d10",-- -2095
x"f7950",-- -2155
x"f4980",-- -2920
x"f2e60",-- -3354
x"f06b0",-- -3989
x"eb6f0",-- -5265
x"e51d0",-- -6883
x"df370",-- -8393
x"de380",-- -8648
x"e1ea0",-- -7702
x"e9810",-- -5759
x"f0710",-- -3983
x"f36f0",-- -3217
x"f2c30",-- -3389
x"f34a0",-- -3254
x"f7f90",-- -2055
x"f94a0",-- -1718
x"fb680",-- -1176
x"023c0",-- 572
x"09c70",-- 2503
x"11650",-- 4453
x"16410",-- 5697
x"164a0",-- 5706
x"118f0",-- 4495
x"0d1d0",-- 3357
x"0b300",-- 2864
x"09880",-- 2440
x"09080",-- 2312
x"078f0",-- 1935
x"05760",-- 1398
x"04b40",-- 1204
x"02440",-- 580
x"fb450",-- -1211
x"f32e0",-- -3282
x"ed830",-- -4733
x"ea240",-- -5596
x"ea8d0",-- -5491
x"ec050",-- -5115
x"ec510",-- -5039
x"eb480",-- -5304
x"ea0a0",-- -5622
x"e9f10",-- -5647
x"e9fc0",-- -5636
x"ea0a0",-- -5622
x"eb880",-- -5240
x"ef8b0",-- -4213
x"f6390",-- -2503
x"fbba0",-- -1094
x"ff9c0",-- -100
x"038b0",-- 907
x"05590",-- 1369
x"07e20",-- 2018
x"0a9b0",-- 2715
x"0d420",-- 3394
x"10160",-- 4118
x"11130",-- 4371
x"12640",-- 4708
x"13720",-- 4978
x"12b30",-- 4787
x"0ef00",-- 3824
x"0a750",-- 2677
x"08c20",-- 2242
x"07830",-- 1923
x"05c70",-- 1479
x"03470",-- 839
x"00960",-- 150
x"fd6f0",-- -657
x"fa410",-- -1471
x"f7fd0",-- -2051
x"f4e10",-- -2847
x"f2e80",-- -3352
x"f16b0",-- -3733
x"f23a0",-- -3526
x"f4570",-- -2985
x"f4d20",-- -2862
x"f54f0",-- -2737
x"f5700",-- -2704
x"f7450",-- -2235
x"f9990",-- -1639
x"fc6b0",-- -917
x"fefa0",-- -262
x"00d50",-- 213
x"03d30",-- 979
x"06f20",-- 1778
x"09ce0",-- 2510
x"0aaa0",-- 2730
x"0af70",-- 2807
x"0bcb0",-- 3019
x"0db00",-- 3504
x"0fa10",-- 4001
x"109b0",-- 4251
x"11300",-- 4400
x"10de0",-- 4318
x"10ca0",-- 4298
x"10c20",-- 4290
x"11290",-- 4393
x"10070",-- 4103
x"0ef70",-- 3831
x"0ea40",-- 3748
x"106b0",-- 4203
x"12f70",-- 4855
x"138a0",-- 5002
x"136a0",-- 4970
x"12370",-- 4663
x"12eb0",-- 4843
x"11e70",-- 4583
x"0c540",-- 3156
x"04430",-- 1091
x"fc4d0",-- -947
x"fa070",-- -1529
x"fc7d0",-- -899
x"fdfb0",-- -517
x"fc050",-- -1019
x"f6610",-- -2463
x"f28a0",-- -3446
x"f06e0",-- -3986
x"ece60",-- -4890
x"e7ca0",-- -6198
x"e2150",-- -7659
x"e1de0",-- -7714
x"e5d10",-- -6703
x"ea290",-- -5591
x"ed240",-- -4828
x"ed430",-- -4797
x"ec5f0",-- -5025
x"ed130",-- -4845
x"f1720",-- -3726
x"f5dd0",-- -2595
x"f9340",-- -1740
x"fdc10",-- -575
x"04910",-- 1169
x"0b880",-- 2952
x"0f030",-- 3843
x"0ec30",-- 3779
x"0c7a0",-- 3194
x"0b300",-- 2864
x"0bdf0",-- 3039
x"0d3a0",-- 3386
x"0de20",-- 3554
x"0cb30",-- 3251
x"0acc0",-- 2764
x"09510",-- 2385
x"07350",-- 1845
x"02940",-- 660
x"fc820",-- -894
x"f7880",-- -2168
x"f5740",-- -2700
x"f5950",-- -2667
x"f4a00",-- -2912
x"f2460",-- -3514
x"eebe0",-- -4418
x"ebe80",-- -5144
x"eab90",-- -5447
x"ea510",-- -5551
x"eaaf0",-- -5457
x"eb450",-- -5307
x"ee320",-- -4558
x"f2060",-- -3578
x"f5160",-- -2794
x"f66c0",-- -2452
x"f8160",-- -2026
x"fb130",-- -1261
x"fea00",-- -352
x"02a00",-- 672
x"05d60",-- 1494
x"09bf0",-- 2495
x"0bc90",-- 3017
x"0cd60",-- 3286
x"0dda0",-- 3546
x"0dd80",-- 3544
x"0d470",-- 3399
x"0bd80",-- 3032
x"0c0f0",-- 3087
x"0ca40",-- 3236
x"0c660",-- 3174
x"0acc0",-- 2764
x"08530",-- 2131
x"05720",-- 1394
x"022f0",-- 559
x"ffdb0",-- -37
x"fd9a0",-- -614
x"fc580",-- -936
x"facd0",-- -1331
x"fa080",-- -1528
x"f9ce0",-- -1586
x"f88c0",-- -1908
x"f7660",-- -2202
x"f6530",-- -2477
x"f6a20",-- -2398
x"f7c60",-- -2106
x"f9770",-- -1673
x"fb6f0",-- -1169
x"fd200",-- -736
x"fec50",-- -315
x"000c0",-- 12
x"01b20",-- 434
x"02ed0",-- 749
x"04410",-- 1089
x"056d0",-- 1389
x"07270",-- 1831
x"08f70",-- 2295
x"09b20",-- 2482
x"0a000",-- 2560
x"09c70",-- 2503
x"099a0",-- 2458
x"093f0",-- 2367
x"09040",-- 2308
x"092b0",-- 2347
x"092b0",-- 2347
x"09290",-- 2345
x"09090",-- 2313
x"08f40",-- 2292
x"091a0",-- 2330
x"08cd0",-- 2253
x"099a0",-- 2458
x"09da0",-- 2522
x"0a7a0",-- 2682
x"0b220",-- 2850
x"0b950",-- 2965
x"0ae50",-- 2789
x"08030",-- 2051
x"06500",-- 1616
x"05830",-- 1411
x"069f0",-- 1695
x"06c80",-- 1736
x"06a90",-- 1705
x"06020",-- 1538
x"04820",-- 1154
x"03330",-- 819
x"004b0",-- 75
x"fd590",-- -679
x"f91a0",-- -1766
x"f6690",-- -2455
x"f5740",-- -2700
x"f5040",-- -2812
x"f4cd0",-- -2867
x"f3d80",-- -3112
x"f3330",-- -3277
x"f1ac0",-- -3668
x"f1110",-- -3823
x"f0f30",-- -3853
x"f1360",-- -3786
x"f2030",-- -3581
x"f3890",-- -3191
x"f6620",-- -2462
x"f8910",-- -1903
x"fa110",-- -1519
x"fa710",-- -1423
x"faad0",-- -1363
x"fb110",-- -1263
x"fb740",-- -1164
x"fc620",-- -926
x"fd880",-- -632
x"feeb0",-- -277
x"00080",-- 8
x"00e30",-- 227
x"01030",-- 259
x"00530",-- 83
x"ff2c0",-- -212
x"fde20",-- -542
x"fd070",-- -761
x"fc620",-- -926
x"fc3f0",-- -961
x"fc6b0",-- -917
x"fcd50",-- -811
x"fd180",-- -744
x"fcd90",-- -807
x"fcc60",-- -826
x"fcaf0",-- -849
x"fcf30",-- -781
x"fd8f0",-- -625
x"fec60",-- -314
x"002b0",-- 43
x"016d0",-- 365
x"027f0",-- 639
x"03420",-- 834
x"04030",-- 1027
x"04340",-- 1076
x"046c0",-- 1132
x"04870",-- 1159
x"04fc0",-- 1276
x"05950",-- 1429
x"05d10",-- 1489
x"05e40",-- 1508
x"05580",-- 1368
x"04bb0",-- 1211
x"03e70",-- 999
x"02fe0",-- 766
x"02190",-- 537
x"016a0",-- 362
x"00c80",-- 200
x"00550",-- 85
x"ffdd0",-- -35
x"ff100",-- -240
x"fe2a0",-- -470
x"fd4a0",-- -694
x"fcaa0",-- -854
x"fc460",-- -954
x"fc250",-- -987
x"fc260",-- -986
x"fc460",-- -954
x"fc690",-- -919
x"fc960",-- -874
x"fc910",-- -879
x"fcaf0",-- -849
x"fccb0",-- -821
x"fd060",-- -762
x"fd950",-- -619
x"fe2f0",-- -465
x"fec50",-- -315
x"ff260",-- -218
x"ff530",-- -173
x"ff3a0",-- -198
x"ff300",-- -208
x"ff2e0",-- -210
x"ff290",-- -215
x"ff510",-- -175
x"ff630",-- -157
x"ff9f0",-- -97
x"ffc20",-- -62
x"ffd60",-- -42
x"ffbc0",-- -68
x"ff850",-- -123
x"ff880",-- -120
x"ff9f0",-- -97
x"00030",-- 3
x"00990",-- 153
x"01490",-- 329
x"01e00",-- 480
x"02890",-- 649
x"03260",-- 806
x"03b50",-- 949
x"04700",-- 1136
x"05350",-- 1333
x"06300",-- 1584
x"073b0",-- 1851
x"086b0",-- 2155
x"09710",-- 2417
x"0a4a0",-- 2634
x"0b040",-- 2820
x"0b990",-- 2969
x"0c250",-- 3109
x"0c980",-- 3224
x"0cde0",-- 3294
x"0cd90",-- 3289
x"0cb80",-- 3256
x"0c270",-- 3111
x"0b620",-- 2914
x"0a6b0",-- 2667
x"091f0",-- 2335
x"07c20",-- 1986
x"06520",-- 1618
x"04ef0",-- 1263
x"03a60",-- 934
x"02500",-- 592
x"01090",-- 265
x"ffd10",-- -47
x"feb70",-- -329
x"fdb50",-- -587
x"fcb10",-- -847
x"fbf80",-- -1032
x"fb4d0",-- -1203
x"faca0",-- -1334
x"fa5d0",-- -1443
x"f9fb0",-- -1541
x"f9ad0",-- -1619
x"f93b0",-- -1733
x"f8de0",-- -1826
x"f87a0",-- -1926
x"f8190",-- -2023
x"f7860",-- -2170
x"f7100",-- -2288
x"f68a0",-- -2422
x"f6030",-- -2557
x"f5980",-- -2664
x"f5570",-- -2729
x"f5330",-- -2765
x"f4fd0",-- -2819
x"f50e0",-- -2802
x"f5270",-- -2777
x"f5750",-- -2699
x"f5bb0",-- -2629
x"f62f0",-- -2513
x"f6cd0",-- -2355
x"f7830",-- -2173
x"f8550",-- -1963
x"f9240",-- -1756
x"f9f80",-- -1544
x"fab20",-- -1358
x"fb7e0",-- -1154
x"fc460",-- -954
x"fd330",-- -717
x"fe080",-- -504
x"febe0",-- -322
x"ff8d0",-- -115
x"00410",-- 65
x"00ca0",-- 202
x"01180",-- 280
x"016a0",-- 362
x"01b20",-- 434
x"02000",-- 512
x"02520",-- 594
x"02820",-- 642
x"02b60",-- 694
x"02e50",-- 741
x"031a0",-- 794
x"035e0",-- 862
x"03720",-- 882
x"03800",-- 896
x"03ad0",-- 941
x"03fe0",-- 1022
x"04350",-- 1077
x"04520",-- 1106
x"04620",-- 1122
x"046c0",-- 1132
x"04660",-- 1126
x"04480",-- 1096
x"043c0",-- 1084
x"04140",-- 1044
x"03dd0",-- 989
x"03ae0",-- 942
x"037e0",-- 894
x"03380",-- 824
x"02c10",-- 705
x"023f0",-- 575
x"01db0",-- 475
x"017b0",-- 379
x"01180",-- 280
x"00ad0",-- 173
x"004b0",-- 75
x"fff30",-- -13
x"ffb20",-- -78
x"ff680",-- -152
x"ff150",-- -235
x"fec50",-- -315
x"fe870",-- -377
x"fe840",-- -380
x"feaf0",-- -337
x"fed70",-- -297
x"fef00",-- -272
x"ff1f0",-- -225
x"ff7b0",-- -133
x"ffd30",-- -45
x"00210",-- 33
x"00910",-- 145
x"01260",-- 294
x"01d10",-- 465
x"02aa0",-- 682
x"03940",-- 916
x"04640",-- 1124
x"05270",-- 1319
x"05ef0",-- 1519
x"06bb0",-- 1723
x"07720",-- 1906
x"081c0",-- 2076
x"08a00",-- 2208
x"09030",-- 2307
x"09450",-- 2373
x"094e0",-- 2382
x"08ef0",-- 2287
x"084b0",-- 2123
x"078d0",-- 1933
x"06a20",-- 1698
x"05b20",-- 1458
x"04c30",-- 1219
x"03d50",-- 981
x"02d20",-- 722
x"01da0",-- 474
x"00eb0",-- 235
x"00000",-- 0
x"ff2e0",-- -210
x"fe6c0",-- -404
x"fdd00",-- -560
x"fd600",-- -672
x"fd1b0",-- -741
x"fce90",-- -791
x"fcb70",-- -841
x"fc710",-- -911
x"fc020",-- -1022
x"fba40",-- -1116
x"fb470",-- -1209
x"fad90",-- -1319
x"fa780",-- -1416
x"fa050",-- -1531
x"f9a60",-- -1626
x"f94a0",-- -1718
x"f8e10",-- -1823
x"f8670",-- -1945
x"f7f40",-- -2060
x"f78b0",-- -2165
x"f7330",-- -2253
x"f7100",-- -2288
x"f6f00",-- -2320
x"f6e60",-- -2330
x"f6df0",-- -2337
x"f6f70",-- -2313
x"f73e0",-- -2242
x"f77f0",-- -2177
x"f7e70",-- -2073
x"f8480",-- -1976
x"f8c10",-- -1855
x"f95e0",-- -1698
x"f9ec0",-- -1556
x"fa7f0",-- -1409
x"fb1f0",-- -1249
x"fbc90",-- -1079
x"fc500",-- -944
x"fcde0",-- -802
x"fd4c0",-- -692
x"fdbf0",-- -577
x"fe3c0",-- -452
x"feb70",-- -329
x"ff440",-- -188
x"ffad0",-- -83
x"001e0",-- 30
x"00ad0",-- 173
x"01420",-- 322
x"01d80",-- 472
x"025c0",-- 604
x"02e60",-- 742
x"03620",-- 866
x"03e50",-- 997
x"04580",-- 1112
x"04c00",-- 1216
x"050e0",-- 1294
x"05540",-- 1364
x"057b0",-- 1403
x"058a0",-- 1418
x"05990",-- 1433
x"05880",-- 1416
x"05800",-- 1408
x"055e0",-- 1374
x"053a0",-- 1338
x"05080",-- 1288
x"04d10",-- 1233
x"047b0",-- 1147
x"042b0",-- 1067
x"03dd0",-- 989
x"03920",-- 914
x"03450",-- 837
x"02f70",-- 759
x"02c10",-- 705
x"02780",-- 632
x"023f0",-- 575
x"01fd0",-- 509
x"01ad0",-- 429
x"01670",-- 359
x"01210",-- 289
x"00e60",-- 230
x"00b60",-- 182
x"009e0",-- 158
x"00700",-- 112
x"00460",-- 70
x"00190",-- 25
x"00000",-- 0
x"fffb0",-- -5
x"fffe0",-- -2
x"001b0",-- 27
x"004b0",-- 75
x"00a20",-- 162
x"01010",-- 257
x"01920",-- 402
x"023a0",-- 570
x"02dc0",-- 732
x"038a0",-- 906
x"04440",-- 1092
x"05170",-- 1303
x"05e70",-- 1511
x"06b90",-- 1721
x"075e0",-- 1886
x"07c20",-- 1986
x"07ef0",-- 2031
x"07db0",-- 2011
x"078d0",-- 1933
x"070b0",-- 1803
x"06760",-- 1654
x"05c60",-- 1478
x"04f20",-- 1266
x"040d0",-- 1037
x"03120",-- 786
x"02030",-- 515
x"00e10",-- 225
x"ffd80",-- -40
x"fedf0",-- -289
x"fe1b0",-- -485
x"fd830",-- -637
x"fd160",-- -746
x"fcd00",-- -816
x"fc9b0",-- -869
x"fc6b0",-- -917
x"fc2f0",-- -977
x"fbe90",-- -1047
x"fb9a0",-- -1126
x"fb5e0",-- -1186
x"fb360",-- -1226
x"fb0e0",-- -1266
x"fadc0",-- -1316
x"faa70",-- -1369
x"fa620",-- -1438
x"fa120",-- -1518
x"f9a80",-- -1624
x"f9420",-- -1726
x"f8d40",-- -1836
x"f8670",-- -1945
x"f8200",-- -2016
x"f7db0",-- -2085
x"f7ad0",-- -2131
x"f7830",-- -2173
x"f7600",-- -2208
x"f74a0",-- -2230
x"f74a0",-- -2230
x"f76d0",-- -2195
x"f7b20",-- -2126
x"f80a0",-- -2038
x"f8700",-- -1936
x"f9010",-- -1791
x"f9970",-- -1641
x"fa390",-- -1479
x"fade0",-- -1314
x"fb790",-- -1159
x"fc1c0",-- -996
x"fcbb0",-- -837
x"fd540",-- -684
x"fddf0",-- -545
x"fe580",-- -424
x"fee10",-- -287
x"ff580",-- -168
x"ffc90",-- -55
x"003f0",-- 63
x"00aa0",-- 170
x"01100",-- 272
x"01810",-- 385
x"01f30",-- 499
x"02670",-- 615
x"02cf0",-- 719
x"03360",-- 822
x"039c0",-- 924
x"03ef0",-- 1007
x"04520",-- 1106
x"04980",-- 1176
x"04c30",-- 1219
x"04ea0",-- 1258
x"05090",-- 1289
x"05100",-- 1296
x"05120",-- 1298
x"04fe0",-- 1278
x"04cd0",-- 1229
x"04be0",-- 1214
x"048c0",-- 1164
x"04580",-- 1112
x"04260",-- 1062
x"03f30",-- 1011
x"03c70",-- 967
x"03920",-- 914
x"03650",-- 869
x"03220",-- 802
x"02e30",-- 739
x"02b10",-- 689
x"027d0",-- 637
x"02580",-- 600
x"021e0",-- 542
x"01da0",-- 474
x"01a90",-- 425
x"016f0",-- 367
x"01330",-- 307
x"00f40",-- 244
x"00ac0",-- 172
x"00870",-- 135
x"00730",-- 115
x"00640",-- 100
x"005d0",-- 93
x"005f0",-- 95
x"00800",-- 128
x"00a00",-- 160
x"00d90",-- 217
x"01310",-- 305
x"01b00",-- 432
x"024b0",-- 587
x"02ef0",-- 751
x"03950",-- 917
x"04430",-- 1091
x"04fe0",-- 1278
x"05b80",-- 1464
x"06700",-- 1648
x"06ea0",-- 1770
x"07490",-- 1865
x"07800",-- 1920
x"07830",-- 1923
x"07560",-- 1878
x"06ff0",-- 1791
x"06870",-- 1671
x"05c60",-- 1478
x"04e50",-- 1253
x"03f10",-- 1009
x"02f00",-- 752
x"01db0",-- 475
x"00c50",-- 197
x"ffd10",-- -47
x"fefd0",-- -259
x"fe3e0",-- -450
x"fd9e0",-- -610
x"fd160",-- -746
x"fcb70",-- -841
x"fc750",-- -907
x"fc3f0",-- -961
x"fc190",-- -999
x"fbec0",-- -1044
x"fbb80",-- -1096
x"fb900",-- -1136
x"fb6a0",-- -1174
x"fb3e0",-- -1218
x"fb070",-- -1273
x"fabe0",-- -1346
x"fa710",-- -1423
x"fa230",-- -1501
x"f9c10",-- -1599
x"f96d0",-- -1683
x"f9240",-- -1756
x"f8cd0",-- -1843
x"f8730",-- -1933
x"f8260",-- -2010
x"f7ea0",-- -2070
x"f7bc0",-- -2116
x"f7930",-- -2157
x"f7920",-- -2158
x"f7b80",-- -2120
x"f7e90",-- -2071
x"f8320",-- -1998
x"f8840",-- -1916
x"f8f00",-- -1808
x"f9660",-- -1690
x"f9e50",-- -1563
x"fa8a0",-- -1398
x"fb2e0",-- -1234
x"fbbd0",-- -1091
x"fc4d0",-- -947
x"fce30",-- -797
x"fd6d0",-- -659
x"fdee0",-- -530
x"fe530",-- -429
x"feb90",-- -327
x"ff360",-- -202
x"ff9c0",-- -100
x"00120",-- 18
x"00910",-- 145
x"00f70",-- 247
x"01790",-- 377
x"01f30",-- 499
x"025f0",-- 607
x"02be0",-- 702
x"031d0",-- 797
x"037b0",-- 891
x"03da0",-- 986
x"04300",-- 1072
x"04690",-- 1129
x"049b0",-- 1179
x"04b80",-- 1208
x"04cd0",-- 1229
x"04c70",-- 1223
x"04ca0",-- 1226
x"04be0",-- 1214
x"04960",-- 1174
x"048a0",-- 1162
x"04730",-- 1139
x"044d0",-- 1101
x"042b0",-- 1067
x"03f80",-- 1016
x"03cb0",-- 971
x"03a40",-- 932
x"03790",-- 889
x"03360",-- 822
x"03040",-- 772
x"02c60",-- 710
x"027b0",-- 635
x"023c0",-- 572
x"01f60",-- 502
x"01b00",-- 432
x"01510",-- 337
x"01030",-- 259
x"00ca0",-- 202
x"00980",-- 152
x"005c0",-- 92
x"00250",-- 37
x"000d0",-- 13
x"fffe0",-- -2
x"fff90",-- -7
x"00070",-- 7
x"001e0",-- 30
x"00390",-- 57
x"007a0",-- 122
x"00ca0",-- 202
x"01120",-- 274
x"01a30",-- 419
x"023f0",-- 575
x"02d40",-- 724
x"035e0",-- 862
x"03e70",-- 999
x"04710",-- 1137
x"05170",-- 1303
x"05c40",-- 1476
x"06300",-- 1584
x"06820",-- 1666
x"06aa0",-- 1706
x"06910",-- 1681
x"06480",-- 1608
x"05e50",-- 1509
x"05650",-- 1381
x"04b40",-- 1204
x"03ee0",-- 1006
x"032c0",-- 812
x"025a0",-- 602
x"01650",-- 357
x"006c0",-- 108
x"ff9e0",-- -98
x"fed50",-- -299
x"fe190",-- -487
x"fd990",-- -615
x"fd3d0",-- -707
x"fce90",-- -791
x"fcad0",-- -851
x"fc820",-- -894
x"fc550",-- -939
x"fc1c0",-- -996
x"fbc70",-- -1081
x"fb850",-- -1147
x"fb620",-- -1182
x"fb360",-- -1226
x"fb040",-- -1276
x"fad90",-- -1319
x"fa9d0",-- -1379
x"fa350",-- -1483
x"f9d00",-- -1584
x"f97e0",-- -1666
x"f9330",-- -1741
x"f8ca0",-- -1846
x"f87d0",-- -1923
x"f8580",-- -1960
x"f8320",-- -1998
x"f8230",-- -2013
x"f8160",-- -2026
x"f81e0",-- -2018
x"f83c0",-- -1988
x"f8670",-- -1945
x"f8a50",-- -1883
x"f90e0",-- -1778
x"f9830",-- -1661
x"f9f10",-- -1551
x"fa670",-- -1433
x"fad90",-- -1319
x"fb3e0",-- -1218
x"fb9e0",-- -1122
x"fc170",-- -1001
x"fc910",-- -879
x"fd130",-- -749
x"fda10",-- -607
x"fe1c0",-- -484
x"fea00",-- -352
x"ff0c0",-- -244
x"ff800",-- -128
x"00000",-- 0
x"008e0",-- 142
x"011a0",-- 282
x"01ad0",-- 429
x"02480",-- 584
x"02ca0",-- 714
x"033d0",-- 829
x"03a10",-- 929
x"03e90",-- 1001
x"04350",-- 1077
x"04620",-- 1122
x"04980",-- 1176
x"04e50",-- 1253
x"04f90",-- 1273
x"050e0",-- 1294
x"05120",-- 1298
x"051a0",-- 1306
x"04ef0",-- 1263
x"04db0",-- 1243
x"04b10",-- 1201
x"04bd0",-- 1213
x"04820",-- 1154
x"048a0",-- 1162
x"04370",-- 1079
x"043e0",-- 1086
x"03c40",-- 964
x"03ea0",-- 1002
x"02ca0",-- 714
x"02160",-- 534
x"04e80",-- 1256
x"03090",-- 777
x"019a0",-- 410
x"018a0",-- 394
x"02990",-- 665
x"024b0",-- 587
x"005f0",-- 95
x"00fa0",-- 250
x"00f90",-- 249
x"00ad0",-- 173
x"00440",-- 68
x"004b0",-- 75
x"00980",-- 152
x"002f0",-- 47
x"00250",-- 37
x"00210",-- 33
x"003f0",-- 63
x"00800",-- 128
x"00b60",-- 182
x"01100",-- 272
x"01510",-- 337
x"01ea0",-- 490
x"024b0",-- 587
x"02d20",-- 722
x"033a0",-- 826
x"03a40",-- 932
x"045c0",-- 1116
x"04fc0",-- 1276
x"056a0",-- 1386
x"05b80",-- 1464
x"060a0",-- 1546
x"05e50",-- 1509
x"05bf0",-- 1471
x"054e0",-- 1358
x"05080",-- 1288
x"049b0",-- 1179
x"03db0",-- 987
x"033d0",-- 829
x"02910",-- 657
x"01cc0",-- 460
x"00e80",-- 232
x"00000",-- 0
x"ff530",-- -173
x"fec80",-- -312
x"fe3a0",-- -454
x"fdef0",-- -529
x"fdae0",-- -594
x"fd6f0",-- -657
x"fd1f0",-- -737
x"fced0",-- -787
x"fcd00",-- -816
x"fc620",-- -926
x"fc230",-- -989
x"fc080",-- -1016
x"fbe50",-- -1051
x"fbbd0",-- -1091
x"fb900",-- -1136
x"fb4c0",-- -1204
x"faf20",-- -1294
x"fa9d0",-- -1379
x"fa4e0",-- -1458
x"fa050",-- -1531
x"f9b70",-- -1609
x"f97a0",-- -1670
x"f95b0",-- -1701
x"f9420",-- -1726
x"f9160",-- -1770
x"f8f70",-- -1801
x"f8eb0",-- -1813
x"f8e80",-- -1816
x"f9290",-- -1751
x"f9590",-- -1703
x"f9b20",-- -1614
x"fa080",-- -1528
x"fa4b0",-- -1461
x"faad0",-- -1363
x"fafc0",-- -1284
x"fb480",-- -1208
x"fba40",-- -1116
x"fc280",-- -984
x"fc8e0",-- -882
x"fd160",-- -746
x"fd860",-- -634
x"fe080",-- -504
x"fe750",-- -395
x"fed70",-- -297
x"ff5d0",-- -163
x"ffd60",-- -42
x"00670",-- 103
x"00e30",-- 227
x"01770",-- 375
x"01fe0",-- 510
x"026b0",-- 619
x"02db0",-- 731
x"031a0",-- 794
x"037b0",-- 891
x"03bd0",-- 957
x"03f90",-- 1017
x"04480",-- 1096
x"04800",-- 1152
x"049e0",-- 1182
x"04b10",-- 1201
x"04b80",-- 1208
x"04a20",-- 1186
x"049b0",-- 1179
x"04760",-- 1142
x"04780",-- 1144
x"04660",-- 1126
x"04460",-- 1094
x"042a0",-- 1066
x"03fb0",-- 1019
x"03d00",-- 976
x"038f0",-- 911
x"03670",-- 871
x"03300",-- 816
x"02fe0",-- 766
x"02cd0",-- 717
x"02890",-- 649
x"024b0",-- 587
x"02000",-- 512
x"01c20",-- 450
x"01680",-- 360
x"011f0",-- 287
x"00df0",-- 223
x"008f0",-- 143
x"00800",-- 128
x"00440",-- 68
x"001e0",-- 30
x"fffb0",-- -5
x"ffdb0",-- -37
x"ffce0",-- -50
x"ffbf0",-- -65
x"ffe40",-- -28
x"ffee0",-- -18
x"fffe0",-- -2
x"00250",-- 37
x"00610",-- 97
x"009d0",-- 157
x"00e40",-- 228
x"014c0",-- 332
x"01bd0",-- 445
x"023c0",-- 572
x"029d0",-- 669
x"03290",-- 809
x"03a80",-- 936
x"043c0",-- 1084
x"04b80",-- 1208
x"04fe0",-- 1278
x"05400",-- 1344
x"053d0",-- 1341
x"053d0",-- 1341
x"04f00",-- 1264
x"04cd0",-- 1229
x"047d0",-- 1149
x"03c10",-- 961
x"03490",-- 841
x"02980",-- 664
x"01df0",-- 479
x"01310",-- 305
x"00700",-- 112
x"ffda0",-- -38
x"ff4c0",-- -180
x"feb60",-- -330
x"fe5a0",-- -422
x"fe070",-- -505
x"fdb30",-- -589
x"fd850",-- -635
x"fd270",-- -729
x"fd010",-- -767
x"fcc60",-- -826
x"fc850",-- -891
x"fc430",-- -957
x"fc120",-- -1006
x"fbea0",-- -1046
x"fba90",-- -1111
x"fb740",-- -1164
x"fb360",-- -1226
x"fae40",-- -1308
x"fa910",-- -1391
x"fa550",-- -1451
x"fa210",-- -1503
x"f9f40",-- -1548
x"f9ab0",-- -1621
x"f98d0",-- -1651
x"f9570",-- -1705
x"f9470",-- -1721
x"f9480",-- -1720
x"f9330",-- -1741
x"f9290",-- -1751
x"f9450",-- -1723
x"f98a0",-- -1654
x"f9bf0",-- -1601
x"fa080",-- -1528
x"fa480",-- -1464
x"faa00",-- -1376
x"faee0",-- -1298
x"fb570",-- -1193
x"fbd60",-- -1066
x"fc350",-- -971
x"fcbe0",-- -834
x"fd3d0",-- -707
x"fdce0",-- -562
x"fe610",-- -415
x"fedc0",-- -292
x"ff670",-- -153
x"ffea0",-- -22
x"00660",-- 102
x"00e10",-- 225
x"01710",-- 369
x"01ef0",-- 495
x"02460",-- 582
x"029e0",-- 670
x"02f40",-- 756
x"034a0",-- 842
x"03900",-- 912
x"03c10",-- 961
x"04000",-- 1024
x"04340",-- 1076
x"044b0",-- 1099
x"046b0",-- 1131
x"04780",-- 1144
x"047b0",-- 1147
x"04890",-- 1161
x"047b0",-- 1147
x"04700",-- 1136
x"04530",-- 1107
x"042b0",-- 1067
x"04200",-- 1056
x"03fd0",-- 1021
x"03c90",-- 969
x"03990",-- 921
x"03670",-- 871
x"03330",-- 819
x"02f70",-- 759
x"02bb0",-- 699
x"02730",-- 627
x"02210",-- 545
x"01da0",-- 474
x"019a0",-- 410
x"01650",-- 357
x"01260",-- 294
x"00ed0",-- 237
x"00b60",-- 182
x"00840",-- 132
x"005f0",-- 95
x"00390",-- 57
x"00230",-- 35
x"001c0",-- 28
x"00030",-- 3
x"fffb0",-- -5
x"00000",-- 0
x"00110",-- 17
x"002d0",-- 45
x"00530",-- 83
x"00800",-- 128
x"00b20",-- 178
x"00ef0",-- 239
x"013f0",-- 319
x"01bd0",-- 445
x"02120",-- 530
x"027d0",-- 637
x"02de0",-- 734
x"034f0",-- 847
x"03ee0",-- 1006
x"04530",-- 1107
x"04ae0",-- 1198
x"04d20",-- 1234
x"04e30",-- 1251
x"04dc0",-- 1244
x"04a70",-- 1191
x"04850",-- 1157
x"04230",-- 1059
x"03c10",-- 961
x"03450",-- 837
x"02ad0",-- 685
x"02190",-- 537
x"016a0",-- 362
x"00cf0",-- 207
x"002f0",-- 47
x"ffbc0",-- -68
x"ff3b0",-- -197
x"fed50",-- -299
x"fe8c0",-- -372
x"fe2d0",-- -467
x"fdec0",-- -532
x"fda80",-- -600
x"fd5d0",-- -675
x"fd110",-- -751
x"fccb0",-- -821
x"fc8e0",-- -882
x"fc550",-- -939
x"fc200",-- -992
x"fbcc0",-- -1076
x"fb9c0",-- -1124
x"fb430",-- -1213
x"faf70",-- -1289
x"faad0",-- -1363
x"fa5c0",-- -1444
x"fa320",-- -1486
x"f9f90",-- -1543
x"f9c20",-- -1598
x"f9940",-- -1644
x"f9750",-- -1675
x"f94d0",-- -1715
x"f93b0",-- -1733
x"f9340",-- -1740
x"f93e0",-- -1730
x"f9570",-- -1705
x"f97a0",-- -1670
x"f9c90",-- -1591
x"fa050",-- -1531
x"fa410",-- -1471
x"fa8e0",-- -1394
x"faeb0",-- -1301
x"fb5b0",-- -1189
x"fbcb0",-- -1077
x"fc480",-- -952
x"fcd00",-- -816
x"fd4f0",-- -689
x"fdd00",-- -560
x"fe570",-- -425
x"fecb0",-- -309
x"ff4e0",-- -178
x"ffd10",-- -47
x"00530",-- 83
x"00c80",-- 200
x"01510",-- 337
x"01c20",-- 450
x"022a0",-- 554
x"02910",-- 657
x"02d40",-- 724
x"03300",-- 816
x"03760",-- 886
x"03bf0",-- 959
x"03e70",-- 999
x"04170",-- 1047
x"04490",-- 1097
x"04660",-- 1126
x"04660",-- 1126
x"04660",-- 1126
x"04620",-- 1122
x"04660",-- 1126
x"045d0",-- 1117
x"04480",-- 1096
x"04300",-- 1072
x"040a0",-- 1034
x"03e40",-- 996
x"03a30",-- 931
x"036c0",-- 876
x"03350",-- 821
x"02fc0",-- 764
x"02ca0",-- 714
x"029d0",-- 669
x"025f0",-- 607
x"02170",-- 535
x"01d00",-- 464
x"01940",-- 404
x"015d0",-- 349
x"011f0",-- 287
x"00e80",-- 232
x"00bb0",-- 187
x"00910",-- 145
x"00640",-- 100
x"00500",-- 80
x"002a0",-- 42
x"00120",-- 18
x"00000",-- 0
x"fff40",-- -12
x"fff90",-- -7
x"00000",-- 0
x"00200",-- 32
x"003f0",-- 63
x"005d0",-- 93
x"008a0",-- 138
x"00b90",-- 185
x"01130",-- 275
x"01650",-- 357
x"01c20",-- 450
x"022b0",-- 555
x"02870",-- 647
x"02ed0",-- 749
x"035d0",-- 861
x"03c60",-- 966
x"040a0",-- 1034
x"044d0",-- 1101
x"04640",-- 1124
x"045f0",-- 1119
x"04490",-- 1097
x"04230",-- 1059
x"03ee0",-- 1006
x"039e0",-- 926
x"033d0",-- 829
x"02cd0",-- 717
x"025c0",-- 604
x"01d00",-- 464
x"013b0",-- 315
x"00ac0",-- 172
x"00280",-- 40
x"ffc60",-- -58
x"ff600",-- -160
x"ff150",-- -235
x"fec10",-- -319
x"fe7d0",-- -387
x"fe3a0",-- -454
x"fdee0",-- -530
x"fdb50",-- -587
x"fd6a0",-- -662
x"fd1b0",-- -741
x"fcd70",-- -809
x"fc8e0",-- -882
x"fc390",-- -967
x"fc030",-- -1021
x"fbbd0",-- -1091
x"fb620",-- -1182
x"fb290",-- -1239
x"fae40",-- -1308
x"faa00",-- -1376
x"fa690",-- -1431
x"fa2b0",-- -1493
x"fa0f0",-- -1521
x"f9ea0",-- -1558
x"f9d30",-- -1581
x"f9bf0",-- -1601
x"f9b30",-- -1613
x"f9c10",-- -1599
x"f9cc0",-- -1588
x"f9f40",-- -1548
x"fa200",-- -1504
x"fa530",-- -1453
x"fa850",-- -1403
x"facd0",-- -1331
x"fb250",-- -1243
x"fb760",-- -1162
x"fbcb0",-- -1077
x"fc350",-- -971
x"fcb10",-- -847
x"fd240",-- -732
x"fda80",-- -600
x"fe260",-- -474
x"fea70",-- -345
x"ff220",-- -222
x"ff990",-- -103
x"00160",-- 22
x"008f0",-- 143
x"01030",-- 259
x"01740",-- 372
x"01d60",-- 470
x"02350",-- 565
x"02800",-- 640
x"02c30",-- 707
x"03080",-- 776
x"034f0",-- 847
x"03830",-- 899
x"03b30",-- 947
x"03e40",-- 996
x"03f10",-- 1009
x"04070",-- 1031
x"04190",-- 1049
x"04160",-- 1046
x"04140",-- 1044
x"040a0",-- 1034
x"04020",-- 1026
x"03e70",-- 999
x"03ce0",-- 974
x"03ad0",-- 941
x"037e0",-- 894
x"03530",-- 851
x"030b0",-- 779
x"02d70",-- 727
x"02980",-- 664
x"02610",-- 609
x"02230",-- 547
x"01db0",-- 475
x"01990",-- 409
x"014a0",-- 330
x"01080",-- 264
x"00c80",-- 200
x"00840",-- 132
x"004d0",-- 77
x"00260",-- 38
x"00020",-- 2
x"ffe20",-- -30
x"ffbc0",-- -68
x"ff9a0",-- -102
x"ff8a0",-- -118
x"ff760",-- -138
x"ff760",-- -138
x"ff7b0",-- -133
x"ff790",-- -135
x"ff990",-- -103
x"ffb00",-- -80
x"ffce0",-- -50
x"fff60",-- -10
x"00200",-- 32
x"00580",-- 88
x"00960",-- 150
x"00da0",-- 218
x"01180",-- 280
x"016c0",-- 364
x"01d10",-- 465
x"022a0",-- 554
x"027d0",-- 637
x"02c80",-- 712
x"03170",-- 791
x"03760",-- 886
x"03b20",-- 946
x"03d10",-- 977
x"03df0",-- 991
x"03e40",-- 996
x"03d30",-- 979
x"03b30",-- 947
x"03970",-- 919
x"03560",-- 854
x"03030",-- 771
x"02ad0",-- 685
x"02500",-- 592
x"01ef0",-- 495
x"018a0",-- 394
x"011c0",-- 284
x"00b60",-- 182
x"004e0",-- 78
x"fff80",-- -8
x"ffb30",-- -77
x"ff5e0",-- -162
x"ff100",-- -240
x"febe0",-- -322
x"fe6c0",-- -404
x"fe210",-- -479
x"fdc60",-- -570
x"fd6f0",-- -657
x"fd240",-- -732
x"fced0",-- -787
x"fc9b0",-- -869
x"fc530",-- -941
x"fc0c0",-- -1012
x"fbc10",-- -1087
x"fb770",-- -1161
x"fb2f0",-- -1233
x"fb0b0",-- -1269
x"faca0",-- -1334
x"faa00",-- -1376
x"fa8a0",-- -1398
x"fa7d0",-- -1411
x"fa6e0",-- -1426
x"fa690",-- -1431
x"fa750",-- -1419
x"fa870",-- -1401
x"fabc0",-- -1348
x"fae10",-- -1311
x"fb110",-- -1263
x"fb4a0",-- -1206
x"fb880",-- -1144
x"fbdb0",-- -1061
x"fc260",-- -986
x"fc7f0",-- -897
x"fcdf0",-- -801
x"fd420",-- -702
x"fdae0",-- -594
x"fe170",-- -489
x"fe800",-- -384
x"feed0",-- -275
x"ff470",-- -185
x"ffbc0",-- -68
x"00170",-- 23
x"007b0",-- 123
x"00eb0",-- 235
x"013b0",-- 315
x"01970",-- 407
x"01e20",-- 482
x"02280",-- 552
x"025d0",-- 605
x"02a80",-- 680
x"02e80",-- 744
x"03080",-- 776
x"032b0",-- 811
x"03420",-- 834
x"03560",-- 854
x"035e0",-- 862
x"03620",-- 866
x"035b0",-- 859
x"03590",-- 857
x"03490",-- 841
x"033a0",-- 826
x"03290",-- 809
x"030d0",-- 781
x"02e00",-- 736
x"02b40",-- 692
x"028a0",-- 650
x"02580",-- 600
x"02210",-- 545
x"01ec0",-- 492
x"01bd0",-- 445
x"01770",-- 375
x"01330",-- 307
x"00ff0",-- 255
x"00bb0",-- 187
x"00760",-- 118
x"00460",-- 70
x"001b0",-- 27
x"fffb0",-- -5
x"ffcc0",-- -52
x"ff9a0",-- -102
x"ff6d0",-- -147
x"ff4e0",-- -178
x"ff330",-- -205
x"ff1d0",-- -227
x"ff100",-- -240
x"ff040",-- -252
x"ff070",-- -249
x"ff070",-- -249
x"ff100",-- -240
x"ff210",-- -223
x"ff240",-- -220
x"ff440",-- -188
x"ff630",-- -157
x"ff800",-- -128
x"ffb20",-- -78
x"ffda0",-- -38
x"000c0",-- 12
x"003f0",-- 63
x"00750",-- 117
x"00bb0",-- 187
x"00f70",-- 247
x"01350",-- 309
x"01790",-- 377
x"01bc0",-- 444
x"02000",-- 512
x"02440",-- 580
x"02840",-- 644
x"02b90",-- 697
x"02ea0",-- 746
x"03260",-- 806
x"03530",-- 851
x"03760",-- 886
x"03830",-- 899
x"038a0",-- 906
x"037b0",-- 891
x"03560",-- 854
x"033d0",-- 829
x"03060",-- 774
x"02cd0",-- 717
x"02800",-- 640
x"02390",-- 569
x"01e20",-- 482
x"01790",-- 377
x"01150",-- 277
x"00b20",-- 178
x"00520",-- 82
x"fffd0",-- -3
x"ff9c0",-- -100
x"ff510",-- -175
x"ff020",-- -254
x"feaf0",-- -337
x"fe660",-- -410
x"fe140",-- -492
x"fdc60",-- -570
x"fd740",-- -652
x"fd290",-- -727
x"fcdf0",-- -801
x"fcaa0",-- -854
x"fc6c0",-- -916
x"fc340",-- -972
x"fbfd0",-- -1027
x"fbd50",-- -1067
x"fb9e0",-- -1122
x"fb7e0",-- -1154
x"fb6c0",-- -1172
x"fb510",-- -1199
x"fb450",-- -1211
x"fb480",-- -1208
x"fb4c0",-- -1204
x"fb570",-- -1193
x"fb6f0",-- -1169
x"fb8b0",-- -1141
x"fbc40",-- -1084
x"fbec0",-- -1044
x"fc2a0",-- -982
x"fc710",-- -911
x"fcc10",-- -831
x"fd020",-- -766
x"fd450",-- -699
x"fda40",-- -604
x"fe000",-- -512
x"fe610",-- -415
x"feaf0",-- -337
x"ff070",-- -249
x"ff600",-- -160
x"ffbc0",-- -68
x"000d0",-- 13
x"00620",-- 98
x"00aa0",-- 170
x"00fc0",-- 252
x"014a0",-- 330
x"01850",-- 389
x"01d10",-- 465
x"01f90",-- 505
x"02260",-- 550
x"025a0",-- 602
x"02780",-- 632
x"02980",-- 664
x"02b70",-- 695
x"02d20",-- 722
x"02db0",-- 731
x"02db0",-- 731
x"02dc0",-- 732
x"02d40",-- 724
x"02c30",-- 707
x"02ad0",-- 685
x"02980",-- 664
x"027a0",-- 634
x"02620",-- 610
x"023c0",-- 572
x"02030",-- 515
x"01db0",-- 475
x"01a90",-- 425
x"01740",-- 372
x"01420",-- 322
x"01100",-- 272
x"00dc0",-- 220
x"00a80",-- 168
x"00760",-- 118
x"00440",-- 68
x"00140",-- 20
x"fff10",-- -15
x"ffbf0",-- -65
x"ffa10",-- -95
x"ff860",-- -122
x"ff6a0",-- -150
x"ff470",-- -185
x"ff310",-- -207
x"ff260",-- -218
x"ff150",-- -235
x"ff130",-- -237
x"ff150",-- -235
x"ff1f0",-- -225
x"ff330",-- -205
x"ff4a0",-- -182
x"ff5d0",-- -163
x"ff830",-- -125
x"ff9a0",-- -102
x"ffba0",-- -70
x"ffea0",-- -22
x"00050",-- 5
x"00320",-- 50
x"005f0",-- 95
x"008c0",-- 140
x"00c00",-- 192
x"00f00",-- 240
x"01210",-- 289
x"01590",-- 345
x"01900",-- 400
x"01ba0",-- 442
x"01f60",-- 502
x"02230",-- 547
x"023e0",-- 574
x"027b0",-- 635
x"02aa0",-- 682
x"02d20",-- 722
x"02f20",-- 754
x"03010",-- 769
x"03120",-- 786
x"031f0",-- 799
x"031c0",-- 796
x"03060",-- 774
x"02fa0",-- 762
x"02d60",-- 726
x"02a20",-- 674
x"02710",-- 625
x"02320",-- 562
x"01f30",-- 499
x"01a40",-- 420
x"01600",-- 352
x"01080",-- 264
x"00ac0",-- 172
x"00570",-- 87
x"00000",-- 0
x"ffb20",-- -78
x"ff5d0",-- -163
x"ff110",-- -239
x"feca0",-- -310
x"fe7d0",-- -387
x"fe3a0",-- -454
x"fdf60",-- -522
x"fdb20",-- -590
x"fd6f0",-- -657
x"fd3a0",-- -710
x"fd070",-- -761
x"fccb0",-- -821
x"fcaa0",-- -854
x"fc7d0",-- -899
x"fc500",-- -944
x"fc260",-- -986
x"fc0a0",-- -1014
x"fbf40",-- -1036
x"fbee0",-- -1042
x"fbe90",-- -1047
x"fbf10",-- -1039
x"fbfd0",-- -1027
x"fc050",-- -1019
x"fc250",-- -987
x"fc480",-- -952
x"fc640",-- -924
x"fc980",-- -872
x"fcd40",-- -812
x"fd0b0",-- -757
x"fd440",-- -700
x"fd8f0",-- -625
x"fdd80",-- -552
x"fe0d0",-- -499
x"fe570",-- -425
x"fe9e0",-- -354
x"feed0",-- -275
x"ff3b0",-- -197
x"ff8a0",-- -118
x"ffd60",-- -42
x"00120",-- 18
x"00520",-- 82
x"00960",-- 150
x"00d20",-- 210
x"01130",-- 275
x"01560",-- 342
x"01810",-- 385
x"01ad0",-- 429
x"01db0",-- 475
x"01f60",-- 502
x"02170",-- 535
x"022f0",-- 559
x"02430",-- 579
x"02580",-- 600
x"025d0",-- 605
x"02620",-- 610
x"025c0",-- 604
x"025a0",-- 602
x"024b0",-- 587
x"02320",-- 562
x"02250",-- 549
x"02070",-- 519
x"01e70",-- 487
x"01bf0",-- 447
x"019a0",-- 410
x"01740",-- 372
x"01490",-- 329
x"01210",-- 289
x"00f50",-- 245
x"00da0",-- 218
x"00b10",-- 177
x"008c0",-- 140
x"006c0",-- 108
x"00430",-- 67
x"00250",-- 37
x"fffb0",-- -5
x"ffdb0",-- -37
x"ffc10",-- -63
x"ffa90",-- -87
x"ff950",-- -107
x"ff8f0",-- -113
x"ff830",-- -125
x"ff6f0",-- -145
x"ff710",-- -143
x"ff710",-- -143
x"ff6c0",-- -148
x"ff760",-- -138
x"ff860",-- -122
x"ff9e0",-- -98
x"ffa90",-- -87
x"ffc10",-- -63
x"ffe50",-- -27
x"fffe0",-- -2
x"00170",-- 23
x"00370",-- 55
x"005d0",-- 93
x"007d0",-- 125
x"009d0",-- 157
x"00c00",-- 192
x"00e10",-- 225
x"00ff0",-- 255
x"01260",-- 294
x"01490",-- 329
x"01710",-- 369
x"01970",-- 407
x"01bf0",-- 447
x"01d60",-- 470
x"01fd0",-- 509
x"02140",-- 532
x"022a0",-- 554
x"023e0",-- 574
x"02410",-- 577
x"024e0",-- 590
x"02460",-- 582
x"02430",-- 579
x"022f0",-- 559
x"02190",-- 537
x"01f40",-- 500
x"01cb0",-- 459
x"019e0",-- 414
x"016d0",-- 365
x"013b0",-- 315
x"00fc0",-- 252
x"00c00",-- 192
x"007f0",-- 127
x"003f0",-- 63
x"fff90",-- -7
x"ffb50",-- -75
x"ff6a0",-- -150
x"ff2b0",-- -213
x"fee40",-- -284
x"fe990",-- -359
x"fe610",-- -415
x"fe1e0",-- -482
x"fde20",-- -542
x"fda40",-- -604
x"fd6f0",-- -657
x"fd340",-- -716
x"fd020",-- -766
x"fcde0",-- -802
x"fcac0",-- -852
x"fc890",-- -887
x"fc670",-- -921
x"fc520",-- -942
x"fc430",-- -957
x"fc2f0",-- -977
x"fc2d0",-- -979
x"fc2f0",-- -977
x"fc410",-- -959
x"fc520",-- -942
x"fc640",-- -924
x"fc820",-- -894
x"fc9e0",-- -866
x"fccf0",-- -817
x"fd060",-- -762
x"fd330",-- -717
x"fd680",-- -664
x"fdae0",-- -594
x"fdea0",-- -534
x"fe1e0",-- -482
x"fe550",-- -427
x"fea20",-- -350
x"fee10",-- -287
x"ff1f0",-- -225
x"ff680",-- -152
x"ffb20",-- -78
x"fff60",-- -10
x"002f0",-- 47
x"00730",-- 115
x"00ac0",-- 172
x"00f50",-- 245
x"01270",-- 295
x"015d0",-- 349
x"018b0",-- 395
x"01ab0",-- 427
x"01d30",-- 467
x"01f80",-- 504
x"02190",-- 537
x"02340",-- 564
x"02490",-- 585
x"024d0",-- 589
x"02580",-- 600
x"025a0",-- 602
x"02620",-- 610
x"02580",-- 600
x"02520",-- 594
x"02430",-- 579
x"022a0",-- 554
x"021c0",-- 540
x"02000",-- 512
x"01ec0",-- 492
x"01d30",-- 467
x"01ba0",-- 442
x"01990",-- 409
x"017b0",-- 379
x"01540",-- 340
x"013d0",-- 317
x"01220",-- 290
x"01030",-- 259
x"00eb0",-- 235
x"00c10",-- 193
x"00a80",-- 168
x"00890",-- 137
x"00700",-- 112
x"00580",-- 88
x"00430",-- 67
x"00280",-- 40
x"00200",-- 32
x"00170",-- 23
x"00140",-- 20
x"001b0",-- 27
x"000f0",-- 15
x"00160",-- 22
x"00190",-- 25
x"00230",-- 35
x"00230",-- 35
x"00280",-- 40
x"00410",-- 65
x"00440",-- 68
x"005d0",-- 93
x"00660",-- 102
x"007d0",-- 125
x"008f0",-- 143
x"00a30",-- 163
x"00bc0",-- 188
x"00cd0",-- 205
x"00d50",-- 213
x"00e30",-- 227
x"01030",-- 259
x"01150",-- 277
x"01270",-- 295
x"013f0",-- 319
x"01510",-- 337
x"01540",-- 340
x"015d0",-- 349
x"01630",-- 355
x"01630",-- 355
x"01590",-- 345
x"01580",-- 344
x"01440",-- 324
x"013b0",-- 315
x"01270",-- 295
x"01090",-- 265
x"00de0",-- 222
x"00af0",-- 175
x"008c0",-- 140
x"00500",-- 80
x"001c0",-- 28
x"fff30",-- -13
x"ffb80",-- -72
x"ff860",-- -122
x"ff510",-- -175
x"ff1a0",-- -230
x"feee0",-- -274
x"feb70",-- -329
x"fe870",-- -377
x"fe530",-- -429
x"fe1c0",-- -484
x"fdee0",-- -530
x"fdbd0",-- -579
x"fd970",-- -617
x"fd720",-- -654
x"fd4e0",-- -690
x"fd310",-- -719
x"fd100",-- -752
x"fcf30",-- -781
x"fcdf0",-- -801
x"fcd00",-- -816
x"fcc00",-- -832
x"fcb90",-- -839
x"fcc10",-- -831
x"fccb0",-- -821
x"fccd0",-- -819
x"fcdf0",-- -801
x"fcf50",-- -779
x"fd0e0",-- -754
x"fd330",-- -717
x"fd560",-- -682
x"fd880",-- -632
x"fdb70",-- -585
x"fddf0",-- -545
x"fe110",-- -495
x"fe4e0",-- -434
x"fe820",-- -382
x"fec10",-- -319
x"fefa0",-- -262
x"ff310",-- -207
x"ff670",-- -153
x"ff9e0",-- -98
x"ffd60",-- -42
x"00050",-- 5
x"00480",-- 72
x"00840",-- 132
x"00bc0",-- 188
x"00de0",-- 222
x"010d0",-- 269
x"01360",-- 310
x"01590",-- 345
x"017e0",-- 382
x"01a40",-- 420
x"01c10",-- 449
x"01df0",-- 479
x"01ef0",-- 495
x"01fb0",-- 507
x"020c0",-- 524
x"020a0",-- 522
x"02070",-- 519
x"01f60",-- 502
x"01ef0",-- 495
x"01df0",-- 479
x"01d10",-- 465
x"01d30",-- 467
x"01bc0",-- 444
x"01b30",-- 435
x"01b20",-- 434
x"018f0",-- 399
x"01740",-- 372
x"015b0",-- 347
x"013f0",-- 319
x"011f0",-- 287
x"01060",-- 262
x"00eb0",-- 235
x"00d90",-- 217
x"00c50",-- 197
x"00ac0",-- 172
x"00930",-- 147
x"006b0",-- 107
x"00580",-- 88
x"00480",-- 72
x"00210",-- 33
x"001e0",-- 30
x"00170",-- 23
x"00070",-- 7
x"00020",-- 2
x"fff80",-- -8
x"00000",-- 0
x"00000",-- 0
x"fffe0",-- -2
x"fffb0",-- -5
x"00140",-- 20
x"00260",-- 38
x"002b0",-- 43
x"00370",-- 55
x"00520",-- 82
x"00620",-- 98
x"006b0",-- 107
x"008c0",-- 140
x"009d0",-- 157
x"00b40",-- 180
x"00be0",-- 190
x"00cb0",-- 203
x"00de0",-- 222
x"00f40",-- 244
x"01030",-- 259
x"01150",-- 277
x"012c0",-- 300
x"01310",-- 305
x"01350",-- 309
x"013a0",-- 314
x"01330",-- 307
x"01350",-- 309
x"012e0",-- 302
x"01180",-- 280
x"01170",-- 279
x"01100",-- 272
x"00fa0",-- 250
x"00eb0",-- 235
x"00d50",-- 213
x"00b10",-- 177
x"00960",-- 150
x"00610",-- 97
x"003e0",-- 62
x"00280",-- 40
x"00000",-- 0
x"ffd60",-- -42
x"ffae0",-- -82
x"ff800",-- -128
x"ff510",-- -175
x"ff350",-- -203
x"ff040",-- -252
x"fee40",-- -284
x"fec00",-- -320
x"fe8e0",-- -370
x"fe660",-- -410
x"fe3e0",-- -450
x"fe140",-- -492
x"fe030",-- -509
x"fde50",-- -539
x"fdc10",-- -575
x"fdab0",-- -597
x"fd920",-- -622
x"fd850",-- -635
x"fd6f0",-- -657
x"fd590",-- -679
x"fd580",-- -680
x"fd560",-- -682
x"fd630",-- -669
x"fd720",-- -654
x"fd810",-- -639
x"fd940",-- -620
x"fda40",-- -604
x"fdc40",-- -572
x"fddd0",-- -547
x"fe000",-- -512
x"fe160",-- -490
x"fe370",-- -457
x"fe690",-- -407
x"fe960",-- -362
x"fec50",-- -315
x"feed0",-- -275
x"ff180",-- -232
x"ff470",-- -185
x"ff740",-- -140
x"ff9c0",-- -100
x"ffc60",-- -58
x"fff30",-- -13
x"000f0",-- 15
x"003e0",-- 62
x"00660",-- 102
x"008a0",-- 138
x"00b20",-- 178
x"00da0",-- 218
x"00f40",-- 244
x"010d0",-- 269
x"01220",-- 290
x"01350",-- 309
x"01510",-- 337
x"01530",-- 339
x"015e0",-- 350
x"01710",-- 369
x"01740",-- 372
x"01770",-- 375
x"017c0",-- 380
x"01770",-- 375
x"016d0",-- 365
x"01650",-- 357
x"01600",-- 352
x"01510",-- 337
x"014e0",-- 334
x"013b0",-- 315
x"01360",-- 310
x"01240",-- 292
x"010d0",-- 269
x"01060",-- 262
x"00f00",-- 240
x"00da0",-- 218
x"00c00",-- 192
x"00bc0",-- 188
x"00a80",-- 168
x"00930",-- 147
x"007d0",-- 125
x"006b0",-- 107
x"005d0",-- 93
x"004b0",-- 75
x"00440",-- 68
x"00430",-- 67
x"002f0",-- 47
x"00320",-- 50
x"00370",-- 55
x"00340",-- 52
x"00350",-- 53
x"003f0",-- 63
x"003e0",-- 62
x"004e0",-- 78
x"005a0",-- 90
x"00610",-- 97
x"00670",-- 103
x"006b0",-- 107
x"007f0",-- 127
x"008a0",-- 138
x"00a00",-- 160
x"00a30",-- 163
x"00b20",-- 178
x"00b90",-- 185
x"00c10",-- 193
x"00dc0",-- 220
x"00e40",-- 228
x"00f40",-- 244
x"01010",-- 257
x"01080",-- 264
x"010d0",-- 269
x"011f0",-- 287
x"01220",-- 290
x"01220",-- 290
x"01210",-- 289
x"01180",-- 280
x"01180",-- 280
x"010d0",-- 269
x"00ff0",-- 255
x"00f90",-- 249
x"00e90",-- 233
x"00e40",-- 228
x"00d70",-- 215
x"00bc0",-- 188
x"00a00",-- 160
x"00870",-- 135
x"00710",-- 113
x"004b0",-- 75
x"001e0",-- 30
x"00000",-- 0
x"ffdf0",-- -33
x"ffb80",-- -72
x"ff990",-- -103
x"ff790",-- -135
x"ff580",-- -168
x"ff330",-- -205
x"ff1c0",-- -228
x"fef50",-- -267
x"fed20",-- -302
x"feb40",-- -332
x"fe980",-- -360
x"fe750",-- -395
x"fe580",-- -424
x"fe410",-- -447
x"fe2f0",-- -465
x"fe1b0",-- -485
x"fe020",-- -510
x"fdf40",-- -524
x"fdec0",-- -532
x"fddb0",-- -549
x"fdd30",-- -557
x"fdd00",-- -560
x"fdda0",-- -550
x"fde90",-- -535
x"fdf60",-- -522
x"fe0c0",-- -500
x"fe0d0",-- -499
x"fe1e0",-- -482
x"fe2f0",-- -465
x"fe3c0",-- -452
x"fe580",-- -424
x"fe7a0",-- -390
x"fe9b0",-- -357
x"febb0",-- -325
x"fed70",-- -297
x"fef50",-- -267
x"ff1a0",-- -230
x"ff3a0",-- -198
x"ff630",-- -157
x"ff8a0",-- -118
x"ffa60",-- -90
x"ffce0",-- -50
x"ffdd0",-- -35
x"fffe0",-- -2
x"00250",-- 37
x"00340",-- 52
x"00530",-- 83
x"00780",-- 120
x"00820",-- 130
x"00980",-- 152
x"00b70",-- 183
x"00c50",-- 197
x"00d40",-- 212
x"00e60",-- 230
x"00f00",-- 240
x"00f70",-- 247
x"01090",-- 265
x"01100",-- 272
x"01080",-- 264
x"01040",-- 260
x"01090",-- 265
x"00ff0",-- 255
x"01010",-- 257
x"01030",-- 259
x"00fc0",-- 252
x"00f50",-- 245
x"00e90",-- 233
x"00e40",-- 228
x"00e10",-- 225
x"00d70",-- 215
x"00c60",-- 198
x"00be0",-- 190
x"00b20",-- 178
x"009e0",-- 158
x"00870",-- 135
x"00760",-- 118
x"00730",-- 115
x"00610",-- 97
x"00640",-- 100
x"00640",-- 100
x"005a0",-- 90
x"005a0",-- 90
x"00570",-- 87
x"00550",-- 85
x"004b0",-- 75
x"00480",-- 72
x"00370",-- 55
x"00430",-- 67
x"00490",-- 73
x"004b0",-- 75
x"00570",-- 87
x"00570",-- 87
x"00530",-- 83
x"00570",-- 87
x"00620",-- 98
x"00730",-- 115
x"00870",-- 135
x"008c0",-- 140
x"00960",-- 150
x"009d0",-- 157
x"00af0",-- 175
x"00be0",-- 190
x"00cb0",-- 203
x"00d20",-- 210
x"00de0",-- 222
x"00d90",-- 217
x"00dc0",-- 220
x"00eb0",-- 235
x"00e90",-- 233
x"00df0",-- 223
x"00d50",-- 213
x"00d90",-- 217
x"00cf0",-- 207
x"00cd0",-- 205
x"00c60",-- 198
x"00c00",-- 192
x"00bc0",-- 188
x"00af0",-- 175
x"009e0",-- 158
x"008c0",-- 140
x"00750",-- 117
x"00580",-- 88
x"00440",-- 68
x"002b0",-- 43
x"000f0",-- 15
x"fff40",-- -12
x"ffdb0",-- -37
x"ffc90",-- -55
x"ffae0",-- -82
x"ff900",-- -112
x"ff6f0",-- -145
x"ff560",-- -170
x"ff3d0",-- -195
x"ff180",-- -232
x"ff0c0",-- -244
x"feff0",-- -257
x"fee40",-- -284
x"fed40",-- -300
x"febe0",-- -322
x"fea00",-- -352
x"fe8f0",-- -369
x"fe820",-- -382
x"fe760",-- -394
x"fe6b0",-- -405
x"fe570",-- -425
x"fe4e0",-- -434
x"fe530",-- -429
x"fe4e0",-- -434
x"fe440",-- -444
x"fe440",-- -444
x"fe410",-- -447
x"fe460",-- -442
x"fe570",-- -425
x"fe5a0",-- -422
x"fe620",-- -414
x"fe780",-- -392
x"fe930",-- -365
x"fead0",-- -339
x"febc0",-- -324
x"fec50",-- -315
x"fee10",-- -287
x"fef70",-- -265
x"ff110",-- -239
x"ff270",-- -217
x"ff310",-- -207
x"ff470",-- -185
x"ff6a0",-- -150
x"ff670",-- -153
x"ff970",-- -105
x"ffe20",-- -30
x"ffad0",-- -83
x"ffe20",-- -30
x"00070",-- 7
x"00070",-- 7
x"002b0",-- 43
x"002d0",-- 45
x"00390",-- 57
x"004e0",-- 78
x"00610",-- 97
x"00700",-- 112
x"00780",-- 120
x"008a0",-- 138
x"009b0",-- 155
x"00990",-- 153
x"00a20",-- 162
x"009d0",-- 157
x"00a30",-- 163
x"00a70",-- 167
x"009d0",-- 157
x"00a20",-- 162
x"008f0",-- 143
x"00990",-- 153
x"00aa0",-- 170
x"008f0",-- 143
x"008c0",-- 140
x"00840",-- 132
x"00760",-- 118
x"007d0",-- 125
x"007d0",-- 125
x"00700",-- 112
x"006b0",-- 107
x"005c0",-- 92
x"005a0",-- 90
x"00500",-- 80
x"00480",-- 72
x"00550",-- 85
x"004e0",-- 78
x"00440",-- 68
x"00490",-- 73
x"004d0",-- 77
x"00430",-- 67
x"00460",-- 70
x"004b0",-- 75
x"00530",-- 83
x"00570",-- 87
x"00580",-- 88
x"005d0",-- 93
x"00640",-- 100
x"00660",-- 102
x"006c0",-- 108
x"007d0",-- 125
x"007d0",-- 125
x"008c0",-- 140
x"00a00",-- 160
x"00a50",-- 165
x"00b70",-- 183
x"00bc0",-- 188
x"00bc0",-- 188
x"00c80",-- 200
x"00cb0",-- 203
x"00c80",-- 200
x"00d40",-- 212
x"00d90",-- 217
x"00d50",-- 213
x"00da0",-- 218
x"00dc0",-- 220
x"00e40",-- 228
x"00e40",-- 228
x"00e10",-- 225
x"00df0",-- 223
x"00e40",-- 228
x"00d90",-- 217
x"00cd0",-- 205
x"00c80",-- 200
x"00bc0",-- 188
x"00a80",-- 168
x"00990",-- 153
x"008f0",-- 143
x"00780",-- 120
x"005d0",-- 93
x"004b0",-- 75
x"003e0",-- 62
x"00230",-- 35
x"000d0",-- 13
x"00020",-- 2
x"fff80",-- -8
x"ffdb0",-- -37
x"ffbd0",-- -67
x"ffa60",-- -90
x"ff950",-- -107
x"ff800",-- -128
x"ff6c0",-- -148
x"ff590",-- -167
x"ff470",-- -185
x"ff380",-- -200
x"ff2b0",-- -213
x"ff1c0",-- -228
x"ff040",-- -252
x"fefd0",-- -259
x"fee80",-- -280
x"fedc0",-- -292
x"fed90",-- -295
x"feca0",-- -310
x"fec60",-- -314
x"febc0",-- -324
x"feb10",-- -335
x"feaa0",-- -342
x"fea80",-- -344
x"fe9e0",-- -354
x"fea50",-- -347
x"febe0",-- -322
x"febb0",-- -325
x"feb70",-- -329
x"feda0",-- -294
x"fede0",-- -290
x"fede0",-- -290
x"fee80",-- -280
x"fef50",-- -267
x"fefd0",-- -259
x"ff020",-- -254
x"ff180",-- -232
x"ff240",-- -220
x"ff2b0",-- -213
x"ff470",-- -185
x"ff5b0",-- -165
x"ff6f0",-- -145
x"ff8a0",-- -118
x"ff990",-- -103
x"ffa60",-- -90
x"ffbc0",-- -68
x"ffd30",-- -45
x"ffd50",-- -43
x"ffe50",-- -27
x"fff60",-- -10
x"00000",-- 0
x"00050",-- 5
x"00070",-- 7
x"00190",-- 25
x"00210",-- 33
x"00280",-- 40
x"00370",-- 55
x"00390",-- 57
x"003e0",-- 62
x"00490",-- 73
x"00520",-- 82
x"005a0",-- 90
x"00520",-- 82
x"00530",-- 83
x"005a0",-- 90
x"00610",-- 97
x"00580",-- 88
x"00570",-- 87
x"005c0",-- 92
x"00530",-- 83
x"005a0",-- 90
x"005d0",-- 93
x"00610",-- 97
x"005f0",-- 95
x"004e0",-- 78
x"004b0",-- 75
x"004e0",-- 78
x"004e0",-- 78
x"00490",-- 73
x"00490",-- 73
x"00440",-- 68
x"004d0",-- 77
x"004e0",-- 78
x"004b0",-- 75
x"00570",-- 87
x"00530",-- 83
x"00610",-- 97
x"00580",-- 88
x"00610",-- 97
x"006b0",-- 107
x"00660",-- 102
x"006b0",-- 107
x"00730",-- 115
x"00760",-- 118
x"007b0",-- 123
x"008e0",-- 142
x"00960",-- 150
x"00990",-- 153
x"00a50",-- 165
x"00b20",-- 178
x"00a20",-- 162
x"00a50",-- 165
x"00b20",-- 178
x"00b20",-- 178
x"00af0",-- 175
x"00b90",-- 185
x"00bb0",-- 187
x"00c00",-- 192
x"00bc0",-- 188
x"00be0",-- 190
x"00b70",-- 183
x"00b90",-- 185
x"00bc0",-- 188
x"00c50",-- 197
x"00b60",-- 182
x"00a80",-- 168
x"00aa0",-- 170
x"009b0",-- 155
x"00a00",-- 160
x"00990",-- 153
x"00960",-- 150
x"008e0",-- 142
x"00870",-- 135
x"00780",-- 120
x"005f0",-- 95
x"00530",-- 83
x"004b0",-- 75
x"003e0",-- 62
x"00280",-- 40
x"00200",-- 32
x"000f0",-- 15
x"fff90",-- -7
x"ffe70",-- -25
x"ffe50",-- -27
x"ffd80",-- -40
x"ffc90",-- -55
x"ffc40",-- -60
x"ffb20",-- -78
x"ffa30",-- -93
x"ff8b0",-- -117
x"ff720",-- -142
x"ff6f0",-- -145
x"ff6c0",-- -148
x"ff5e0",-- -162
x"ff590",-- -167
x"ff4c0",-- -180
x"ff360",-- -202
x"ff2b0",-- -213
x"ff1f0",-- -225
x"ff110",-- -239
x"ff130",-- -237
x"ff0e0",-- -242
x"ff0b0",-- -245
x"ff040",-- -252
x"ff040",-- -252
x"ff070",-- -249
x"ff070",-- -249
x"ff170",-- -233
x"ff150",-- -235
x"ff180",-- -232
x"ff240",-- -220
x"ff2e0",-- -210
x"ff350",-- -203
x"ff310",-- -207
x"ff360",-- -202
x"ff380",-- -200
x"ff490",-- -183
x"ff470",-- -185
x"ff580",-- -168
x"ff680",-- -152
x"ff6d0",-- -147
x"ff880",-- -120
x"ff920",-- -110
x"ffa10",-- -95
x"ffa30",-- -93
x"ffa90",-- -87
x"ffb50",-- -75
x"ffb00",-- -80
x"ffbf0",-- -65
x"ffd60",-- -42
x"ffdf0",-- -33
x"ffe20",-- -30
x"ffea0",-- -22
x"fff60",-- -10
x"fffb0",-- -5
x"fffb0",-- -5
x"00080",-- 8
x"000c0",-- 12
x"00160",-- 22
x"00190",-- 25
x"001b0",-- 27
x"001e0",-- 30
x"001c0",-- 28
x"00250",-- 37
x"00250",-- 37
x"00210",-- 33
x"00280",-- 40
x"00300",-- 48
x"00340",-- 52
x"00410",-- 65
x"00490",-- 73
x"004e0",-- 78
x"00490",-- 73
x"00410",-- 65
x"00460",-- 70
x"004b0",-- 75
x"00480",-- 72
x"004b0",-- 75
x"00520",-- 82
x"00520",-- 82
x"00500",-- 80
x"00530",-- 83
x"00530",-- 83
x"00530",-- 83
x"005a0",-- 90
x"006b0",-- 107
x"006b0",-- 107
x"006e0",-- 110
x"00710",-- 113
x"006c0",-- 108
x"007a0",-- 122
x"007d0",-- 125
x"00760",-- 118
x"007d0",-- 125
x"00840",-- 132
x"00800",-- 128
x"008f0",-- 143
x"00850",-- 133
x"00840",-- 132
x"008f0",-- 143
x"00930",-- 147
x"00930",-- 147
x"008c0",-- 140
x"00960",-- 150
x"00980",-- 152
x"008c0",-- 140
x"00940",-- 148
x"00910",-- 145
x"00870",-- 135
x"008e0",-- 142
x"00960",-- 150
x"00980",-- 152
x"008c0",-- 140
x"007d0",-- 125
x"00840",-- 132
x"008a0",-- 138
x"007b0",-- 123
x"007d0",-- 125
x"00780",-- 120
x"00700",-- 112
x"00700",-- 112
x"006e0",-- 110
x"00640",-- 100
x"00550",-- 85
x"00500",-- 80
x"004b0",-- 75
x"003e0",-- 62
x"00300",-- 48
x"002a0",-- 42
x"00160",-- 22
x"000d0",-- 13
x"00020",-- 2
x"fffd0",-- -3
x"fffe0",-- -2
x"fff30",-- -13
x"ffd80",-- -40
x"ffd50",-- -43
x"ffc20",-- -62
x"ffc10",-- -63
x"ffa90",-- -87
x"ffb50",-- -75
x"ff8a0",-- -118
x"ff990",-- -103
x"ff530",-- -173
x"ff760",-- -138
x"ff220",-- -222
x"ff4e0",-- -178
x"feca0",-- -310
x"ff110",-- -239
x"fe490",-- -439
x"ff010",-- -255
x"fa120",-- -1518
x"eaca0",-- -5430
x"f5100",-- -2800
x"05170",-- 1303
x"00e30",-- 227
x"fe260",-- -474
x"023f0",-- 575
x"00700",-- 112
x"fe9e0",-- -354
x"01cc0",-- 460
x"ff9c0",-- -100
x"ffd10",-- -47
x"fe490",-- -439
x"fdf10",-- -527
x"00dc0",-- 220
x"fecf0",-- -305
x"00660",-- 102
x"04530",-- 1107
x"fea20",-- -350
x"f7220",-- -2270
x"fc700",-- -912
x"00340",-- 52
x"fe960",-- -362
x"ffee0",-- -18
x"fa390",-- -1479
x"f9f30",-- -1549
x"00e40",-- 228
x"fd590",-- -679
x"fc640",-- -924
x"01e70",-- 487
x"00aa0",-- 170
x"ffd80",-- -40
x"009e0",-- 158
x"fe410",-- -447
x"00160",-- 22
x"04120",-- 1042
x"08250",-- 2085
x"08c50",-- 2245
x"04f20",-- 1266
x"017c0",-- 380
x"01bf0",-- 447
x"01290",-- 297
x"01f80",-- 504
x"02e50",-- 741
x"00610",-- 97
x"01360",-- 310
x"03760",-- 886
x"01040",-- 260
x"00dc0",-- 220
x"ff010",-- -255
x"fb9f0",-- -1121
x"fc960",-- -874
x"01880",-- 392
x"02580",-- 600
x"00280",-- 40
x"001c0",-- 28
x"febb0",-- -325
x"ffef0",-- -17
x"00cf0",-- 207
x"00ac0",-- 172
x"02c00",-- 704
x"03650",-- 869
x"014e0",-- 334
x"01f90",-- 505
x"03d30",-- 979
x"021c0",-- 540
x"ff970",-- -105
x"fd490",-- -695
x"fe4d0",-- -435
x"fd8b0",-- -629
x"fc5f0",-- -929
x"fd2e0",-- -722
x"fce40",-- -796
x"fab60",-- -1354
x"fa990",-- -1383
x"fd1d0",-- -739
x"fd790",-- -647
x"febe0",-- -322
x"ff620",-- -158
x"028a0",-- 650
x"03440",-- 836
x"03040",-- 772
x"04320",-- 1074
x"04990",-- 1177
x"05720",-- 1394
x"08210",-- 2081
x"0a6e0",-- 2670
x"0a750",-- 2677
x"09560",-- 2390
x"09a10",-- 2465
x"094a0",-- 2378
x"09080",-- 2312
x"0a460",-- 2630
x"07fd0",-- 2045
x"05d50",-- 1493
x"05b80",-- 1464
x"04320",-- 1074
x"01ef0",-- 495
x"01c10",-- 449
x"ff130",-- -237
x"fc430",-- -957
x"fd090",-- -759
x"fd5b0",-- -677
x"fbc60",-- -1082
x"fa250",-- -1499
x"f9b20",-- -1614
x"f9180",-- -1768
x"f8b40",-- -1868
x"f93e0",-- -1730
x"f9cb0",-- -1589
x"f9160",-- -1770
x"f8bc0",-- -1860
x"f8930",-- -1901
x"f95c0",-- -1700
x"f9fe0",-- -1538
x"f91d0",-- -1763
x"f9900",-- -1648
x"fb200",-- -1248
x"fc3c0",-- -964
x"fc580",-- -936
x"fc7f0",-- -897
x"fd2a0",-- -726
x"fde90",-- -535
x"fe070",-- -505
x"ff0c0",-- -244
x"feca0",-- -310
x"fe140",-- -492
x"fe8c0",-- -372
x"fe820",-- -382
x"ff7b0",-- -133
x"ff1f0",-- -225
x"fe300",-- -464
x"feda0",-- -294
x"fee80",-- -280
x"fe1b0",-- -485
x"fe110",-- -495
x"fe990",-- -359
x"fd470",-- -697
x"fca80",-- -856
x"fcb10",-- -847
x"fda10",-- -607
x"fe0a0",-- -502
x"fcfa0",-- -774
x"fd440",-- -700
x"fec30",-- -317
x"004e0",-- 78
x"00570",-- 87
x"01290",-- 297
x"02b10",-- 689
x"02b40",-- 692
x"04280",-- 1064
x"06820",-- 1666
x"07260",-- 1830
x"06d20",-- 1746
x"066c0",-- 1644
x"07680",-- 1896
x"0ab40",-- 2740
x"0abe0",-- 2750
x"0b3b0",-- 2875
x"0deb0",-- 3563
x"0dd50",-- 3541
x"0d860",-- 3462
x"0e860",-- 3718
x"0fc20",-- 4034
x"10ed0",-- 4333
x"12230",-- 4643
x"115e0",-- 4446
x"12660",-- 4710
x"12590",-- 4697
x"11e20",-- 4578
x"13ad0",-- 5037
x"14370",-- 5175
x"14140",-- 5140
x"15080",-- 5384
x"14c50",-- 5317
x"118a0",-- 4490
x"0b5d0",-- 2909
x"06ca0",-- 1738
x"08080",-- 2056
x"091f0",-- 2335
x"05290",-- 1321
x"00cf0",-- 207
x"fde40",-- -540
x"f9d30",-- -1581
x"f5b10",-- -2639
x"f28c0",-- -3444
x"ee670",-- -4505
x"e9660",-- -5786
x"e66f0",-- -6545
x"e68a0",-- -6518
x"e6f10",-- -6415
x"e3de0",-- -7202
x"df3b0",-- -8389
x"ddae0",-- -8786
x"dfa70",-- -8281
x"e3130",-- -7405
x"e63c0",-- -6596
x"e8730",-- -6029
x"ea3f0",-- -5569
x"ecc60",-- -4922
x"f01c0",-- -4068
x"f5520",-- -2734
x"f8cd0",-- -1843
x"fa2b0",-- -1493
x"fcb60",-- -842
x"00930",-- 147
x"033b0",-- 827
x"034f0",-- 847
x"03800",-- 896
x"03440",-- 836
x"03f90",-- 1017
x"04620",-- 1122
x"04e30",-- 1251
x"039a0",-- 922
x"007a0",-- 122
x"fcd40",-- -812
x"fad50",-- -1323
x"f9df0",-- -1569
x"f6df0",-- -2337
x"f41e0",-- -3042
x"f1e80",-- -3608
x"f0120",-- -4078
x"ee000",-- -4608
x"ec300",-- -5072
x"ebac0",-- -5204
x"eb2e0",-- -5330
x"eb4c0",-- -5300
x"ed700",-- -4752
x"f05f0",-- -4001
x"f1900",-- -3696
x"f2990",-- -3431
x"f5130",-- -2797
x"f8b20",-- -1870
x"fcaa0",-- -854
x"00410",-- 65
x"03a80",-- 936
x"06620",-- 1634
x"08d40",-- 2260
x"0b260",-- 2854
x"0df60",-- 3574
x"10310",-- 4145
x"113f0",-- 4415
x"12660",-- 4710
x"145a0",-- 5210
x"15690",-- 5481
x"148e0",-- 5262
x"13590",-- 4953
x"13030",-- 4867
x"13090",-- 4873
x"130e0",-- 4878
x"12ac0",-- 4780
x"11aa0",-- 4522
x"0fa80",-- 4008
x"0f720",-- 3954
x"10480",-- 4168
x"0fc80",-- 4040
x"0e2c0",-- 3628
x"0d830",-- 3459
x"0f920",-- 3986
x"134f0",-- 4943
x"14f00",-- 5360
x"151d0",-- 5405
x"151f0",-- 5407
x"17a60",-- 6054
x"1c680",-- 7272
x"1e720",-- 7794
x"1db20",-- 7602
x"1b2b0",-- 6955
x"1be20",-- 7138
x"198c0",-- 6540
x"14ae0",-- 5294
x"0db50",-- 3509
x"094a0",-- 2378
x"07da0",-- 2010
x"043c0",-- 1084
x"01710",-- 369
x"fc210",-- -991
x"f4c50",-- -2875
x"eba60",-- -5210
x"e6960",-- -6506
x"e3480",-- -7352
x"de4e0",-- -8626
x"daaa0",-- -9558
x"d8230",-- -10205
x"d7b90",-- -10311
x"d64c0",-- -10676
x"d6780",-- -10632
x"d6c90",-- -10551
x"d8230",-- -10205
x"dc5b0",-- -9125
x"e2710",-- -7567
x"ea820",-- -5502
x"ef6f0",-- -4241
x"f38d0",-- -3187
x"f82a0",-- -2006
x"fe5d0",-- -419
x"04280",-- 1064
x"087d0",-- 2173
x"0cff0",-- 3327
x"0fd50",-- 4053
x"10a20",-- 4258
x"0f650",-- 3941
x"11530",-- 4435
x"11df0",-- 4575
x"0df10",-- 3569
x"0abd0",-- 2749
x"09ad0",-- 2477
x"0a1b0",-- 2587
x"041e0",-- 1054
x"fc3a0",-- -966
x"f5df0",-- -2593
x"f1ef0",-- -3601
x"eec00",-- -4416
x"ec7e0",-- -4994
x"eac30",-- -5437
x"e5cf0",-- -6705
x"e1b00",-- -7760
x"e02d0",-- -8147
x"e1630",-- -7837
x"e1ba0",-- -7750
x"e19d0",-- -7779
x"e4060",-- -7162
x"e8d50",-- -5931
x"eda60",-- -4698
x"f0bc0",-- -3908
x"f4e30",-- -2845
x"f67a0",-- -2438
x"f9bc0",-- -1604
x"00190",-- 25
x"09360",-- 2358
x"0e700",-- 3696
x"0ea40",-- 3748
x"0fff0",-- 4095
x"11f80",-- 4600
x"15220",-- 5410
x"154a0",-- 5450
x"16f70",-- 5879
x"16480",-- 5704
x"155b0",-- 5467
x"135b0",-- 4955
x"125c0",-- 4700
x"0f5e0",-- 3934
x"0b210",-- 2849
x"091f0",-- 2335
x"076d0",-- 1901
x"08580",-- 2136
x"04cf0",-- 1231
x"032b0",-- 811
x"01fd0",-- 509
x"02200",-- 544
x"04910",-- 1169
x"05c70",-- 1479
x"08e50",-- 2277
x"06250",-- 1573
x"08200",-- 2080
x"0ce60",-- 3302
x"14550",-- 5205
x"18db0",-- 6363
x"1a200",-- 6688
x"1dc10",-- 7617
x"210f0",-- 8463
x"28160",-- 10262
x"2ce30",-- 11491
x"31050",-- 12549
x"2ed10",-- 11985
x"2d580",-- 11608
x"2c340",-- 11316
x"28d60",-- 10454
x"21bf0",-- 8639
x"17460",-- 5958
x"0d180",-- 3352
x"04e50",-- 1253
x"02490",-- 585
x"ffad0",-- -83
x"f6350",-- -2507
x"e9630",-- -5789
x"ddd30",-- -8749
x"d8470",-- -10169
x"d26f0",-- -11665
x"ce100",-- -12784
x"c9b10",-- -13903
x"c5d60",-- -14890
x"c5a50",-- -14939
x"c7ff0",-- -14337
x"cae50",-- -13595
x"cba40",-- -13404
x"cf520",-- -12462
x"d5ed0",-- -10771
x"e1ba0",-- -7750
x"ecdf0",-- -4897
x"f5ec0",-- -2580
x"fbb50",-- -1099
x"01cc0",-- 460
x"090e0",-- 2318
x"10430",-- 4163
x"18040",-- 6148
x"1cb90",-- 7353
x"1e7f0",-- 7807
x"1e3b0",-- 7739
x"1da50",-- 7589
x"1b1f0",-- 6943
x"171f0",-- 5919
x"135e0",-- 4958
x"0f590",-- 3929
x"0a960",-- 2710
x"049d0",-- 1181
x"fea50",-- -347
x"f4ca0",-- -2870
x"ebcf0",-- -5169
x"e5d30",-- -6701
x"e2000",-- -7680
x"ddd60",-- -8746
x"d9930",-- -9837
x"d7430",-- -10429
x"d46c0",-- -11156
x"d45d0",-- -11171
x"d5310",-- -10959
x"d8800",-- -10112
x"dcdf0",-- -8993
x"e2300",-- -7632
x"e84c0",-- -6068
x"ee7a0",-- -4486
x"f4f00",-- -2832
x"f96d0",-- -1683
x"ff300",-- -208
x"059e0",-- 1438
x"0dd10",-- 3537
x"14610",-- 5217
x"180c0",-- 6156
x"1aef0",-- 6895
x"1b3f0",-- 6975
x"1cd30",-- 7379
x"1d920",-- 7570
x"1d560",-- 7510
x"1b460",-- 6982
x"18be0",-- 6334
x"16390",-- 5689
x"11800",-- 4480
x"0c7f0",-- 3199
x"06050",-- 1541
x"01900",-- 400
x"fe260",-- -474
x"fc120",-- -1006
x"f9970",-- -1641
x"f7060",-- -2298
x"f59d0",-- -2659
x"f4f80",-- -2824
x"f77f0",-- -2177
x"fa840",-- -1404
x"fef20",-- -270
x"022f0",-- 559
x"07d30",-- 2003
x"0c9d0",-- 3229
x"10130",-- 4115
x"149b0",-- 5275
x"1ae30",-- 6883
x"22bd0",-- 8893
x"28480",-- 10312
x"2ea70",-- 11943
x"33350",-- 13109
x"366b0",-- 13931
x"38010",-- 14337
x"3ace0",-- 15054
x"3b8e0",-- 15246
x"3a100",-- 14864
x"34f60",-- 13558
x"303b0",-- 12347
x"26130",-- 9747
x"16d90",-- 5849
x"06200",-- 1568
x"fb1b0",-- -1253
x"f61b0",-- -2533
x"efc40",-- -4156
x"e97a0",-- -5766
x"dd820",-- -8830
x"d2080",-- -11768
x"c6090",-- -14839
x"c2220",-- -15838
x"c02e0",-- -16338
x"bdb90",-- -16967
x"bcf60",-- -17162
x"c1700",-- -16016
x"c8510",-- -14255
x"cbfa0",-- -13318
x"d1430",-- -11965
x"d87b0",-- -10117
x"e2c80",-- -7480
x"ef660",-- -4250
x"fe930",-- -365
x"0b4f0",-- 2895
x"12f90",-- 4857
x"18570",-- 6231
x"1e000",-- 7680
x"248d0",-- 9357
x"28d60",-- 10454
x"2ab10",-- 10929
x"29de0",-- 10718
x"275f0",-- 10079
x"23240",-- 8996
x"1a310",-- 6705
x"0f6c0",-- 3948
x"05ec0",-- 1516
x"ff740",-- -140
x"f9420",-- -1726
x"f11f0",-- -3809
x"e7770",-- -6281
x"dc9c0",-- -9060
x"d3b40",-- -11340
x"ce400",-- -12736
x"cb000",-- -13568
x"c9d40",-- -13868
x"c8d50",-- -14123
x"caf60",-- -13578
x"cd840",-- -12924
x"d2060",-- -11770
x"d7d10",-- -10287
x"defa0",-- -8454
x"e73b0",-- -6341
x"f0a70",-- -3929
x"fc4d0",-- -947
x"05170",-- 1303
x"0c0a0",-- 3082
x"10c80",-- 4296
x"175f0",-- 5983
x"1c980",-- 7320
x"20ef0",-- 8431
x"24570",-- 9303
x"259e0",-- 9630
x"24600",-- 9312
x"20190",-- 8217
x"1c200",-- 7200
x"167f0",-- 5759
x"11260",-- 4390
x"0c540",-- 3156
x"07ee0",-- 2030
x"02710",-- 625
x"faeb0",-- -1301
x"f44b0",-- -2997
x"ef180",-- -4328
x"ebf20",-- -5134
x"ea650",-- -5531
x"eb070",-- -5369
x"eccf0",-- -4913
x"ee9e0",-- -4450
x"f1e00",-- -3616
x"f6190",-- -2535
x"fc530",-- -941
x"02d60",-- 726
x"0b470",-- 2887
x"150e0",-- 5390
x"1e2f0",-- 7727
x"260c0",-- 9740
x"28920",-- 10386
x"2b970",-- 11159
x"2f550",-- 12117
x"37c80",-- 14280
x"3e470",-- 15943
x"3fb90",-- 16313
x"3d8c0",-- 15756
x"38890",-- 14473
x"397f0",-- 14719
x"39660",-- 14694
x"376e0",-- 14190
x"2cd90",-- 11481
x"21bc0",-- 8636
x"1b5f0",-- 7007
x"11400",-- 4416
x"ffdf0",-- -33
x"e88d0",-- -6003
x"da1f0",-- -9697
x"d5960",-- -10858
x"d9070",-- -9977
x"d6b90",-- -10567
x"cc330",-- -13261
x"c1160",-- -16106
x"bbd50",-- -17451
x"be530",-- -16813
x"c28d0",-- -15731
x"c84a0",-- -14262
x"ccb70",-- -13129
x"d4b40",-- -11084
x"dee90",-- -8471
x"eb920",-- -5230
x"f34a0",-- -3254
x"f80d0",-- -2035
x"018b0",-- 395
x"0f970",-- 3991
x"1f050",-- 7941
x"27f50",-- 10229
x"2aec0",-- 10988
x"29870",-- 10631
x"28570",-- 10327
x"27ad0",-- 10157
x"255f0",-- 9567
x"20110",-- 8209
x"18400",-- 6208
x"0fe40",-- 4068
x"06200",-- 1568
x"fa0f0",-- -1521
x"e9ce0",-- -5682
x"dc5f0",-- -9121
x"d5d60",-- -10794
x"d4b00",-- -11088
x"d28a0",-- -11638
x"cbb60",-- -13386
x"c6dd0",-- -14627
x"c2420",-- -15806
x"c4580",-- -15272
x"c9690",-- -13975
x"d19a0",-- -11878
x"d8940",-- -10092
x"dfa20",-- -8286
x"eaa80",-- -5464
x"f3dd0",-- -3107
x"fb220",-- -1246
x"01db0",-- 475
x"0bad0",-- 2989
x"17150",-- 5909
x"20430",-- 8259
x"22c70",-- 8903
x"25d20",-- 9682
x"219b0",-- 8603
x"200e0",-- 8206
x"1f190",-- 7961
x"1d2d0",-- 7469
x"18a20",-- 6306
x"0dc40",-- 3524
x"07f80",-- 2040
x"02210",-- 545
x"fe2d0",-- -467
x"f2da0",-- -3366
x"e9e70",-- -5657
x"e51d0",-- -6883
x"e5000",-- -6912
x"e6350",-- -6603
x"e5520",-- -6830
x"e5520",-- -6830
x"e3750",-- -7307
x"e7920",-- -6254
x"ef830",-- -4221
x"f8be0",-- -1858
x"ffa30",-- -93
x"05760",-- 1398
x"0e2d0",-- 3629
x"17080",-- 5896
x"1e770",-- 7799
x"24f90",-- 9465
x"2aa40",-- 10916
x"314b0",-- 12619
x"38240",-- 14372
x"3c480",-- 15432
x"3a180",-- 14872
x"33f30",-- 13299
x"30330",-- 12339
x"32830",-- 12931
x"33e40",-- 13284
x"2e2c0",-- 11820
x"25fa0",-- 9722
x"202d0",-- 8237
x"1f440",-- 8004
x"1acd0",-- 6861
x"11860",-- 4486
x"07540",-- 1876
x"01ef0",-- 495
x"01d30",-- 467
x"f91d0",-- -1763
x"e8190",-- -6119
x"d6b50",-- -10571
x"cf820",-- -12414
x"d5a20",-- -10846
x"dce90",-- -8983
x"e1040",-- -7932
x"dbb90",-- -9287
x"d6260",-- -10714
x"d8850",-- -10107
x"de7b0",-- -8581
x"e4290",-- -7127
x"e6b40",-- -6476
x"ed7f0",-- -4737
x"f6910",-- -2415
x"ffe20",-- -30
x"068b0",-- 1675
x"089a0",-- 2202
x"07a90",-- 1961
x"0b760",-- 2934
x"15090",-- 5385
x"1cac0",-- 7340
x"1d760",-- 7542
x"19550",-- 6485
x"163c0",-- 5692
x"11680",-- 4456
x"0b400",-- 2880
x"02410",-- 577
x"f8e10",-- -1823
x"f2ac0",-- -3412
x"ef270",-- -4313
x"e9e70",-- -5657
x"e0870",-- -8057
x"d6920",-- -10606
x"cedc0",-- -12580
x"cd500",-- -12976
x"d2970",-- -11625
x"d9590",-- -9895
x"dbf10",-- -9231
x"dc640",-- -9116
x"df780",-- -8328
x"e4f80",-- -6920
x"ec6c0",-- -5012
x"f3570",-- -3241
x"faac0",-- -1364
x"01cc0",-- 460
x"08db0",-- 2267
x"0eb80",-- 3768
x"11a50",-- 4517
x"11920",-- 4498
x"11990",-- 4505
x"14160",-- 5142
x"16af0",-- 5807
x"16860",-- 5766
x"11800",-- 4480
x"0a660",-- 2662
x"041b0",-- 1051
x"ff4e0",-- -178
x"f8af0",-- -1873
x"f4370",-- -3017
x"f0ca0",-- -3894
x"f0a30",-- -3933
x"eed00",-- -4400
x"eb010",-- -5375
x"e8ad0",-- -5971
x"e6e70",-- -6425
x"ea050",-- -5627
x"ef4c0",-- -4276
x"f6820",-- -2430
x"faad0",-- -1363
x"fd4f0",-- -689
x"01450",-- 325
x"06be0",-- 1726
x"0cff0",-- 3327
x"12e50",-- 4837
x"177b0",-- 6011
x"1c090",-- 7177
x"20950",-- 8341
x"236e0",-- 9070
x"24b10",-- 9393
x"23dd0",-- 9181
x"240a0",-- 9226
x"24a40",-- 9380
x"267e0",-- 9854
x"27030",-- 9987
x"227a0",-- 8826
x"1bee0",-- 7150
x"17130",-- 5907
x"16b60",-- 5814
x"16460",-- 5702
x"13330",-- 4915
x"11900",-- 4496
x"11cd0",-- 4557
x"15d70",-- 5591
x"162a0",-- 5674
x"13600",-- 4960
x"0db30",-- 3507
x"0a280",-- 2600
x"07bc0",-- 1980
x"03090",-- 777
x"fada0",-- -1318
x"ec620",-- -5022
x"e6580",-- -6568
x"e86a0",-- -6038
x"f1810",-- -3711
x"f0f80",-- -3848
x"e8fa0",-- -5894
x"e1b80",-- -7752
x"dff60",-- -8202
x"e5050",-- -6907
x"e70e0",-- -6386
x"e8820",-- -6014
x"e80f0",-- -6129
x"eccb0",-- -4917
x"f37c0",-- -3204
x"fabe0",-- -1346
x"fc140",-- -1004
x"fc8e0",-- -882
x"ffdf0",-- -33
x"06d60",-- 1750
x"0e930",-- 3731
x"10c80",-- 4296
x"10e10",-- 4321
x"0dba0",-- 3514
x"0ca50",-- 3237
x"09df0",-- 2527
x"04910",-- 1169
x"fadc0",-- -1316
x"f3890",-- -3191
x"f1250",-- -3803
x"ef2c0",-- -4308
x"e8cd0",-- -5939
x"df520",-- -8366
x"dae90",-- -9495
x"db570",-- -9385
x"dd750",-- -8843
x"e0260",-- -8154
x"e4620",-- -7070
x"e6440",-- -6588
x"e8580",-- -6056
x"ec2d0",-- -5075
x"f2de0",-- -3362
x"f7100",-- -2288
x"f9f10",-- -1551
x"ff380",-- -200
x"05290",-- 1321
x"09650",-- 2405
x"0b650",-- 2917
x"0bb30",-- 2995
x"0b4c0",-- 2892
x"0bbc0",-- 3004
x"0bdb0",-- 3035
x"0b0e0",-- 2830
x"06fe0",-- 1790
x"022b0",-- 555
x"fd270",-- -729
x"fa710",-- -1423
x"f78e0",-- -2162
x"f4f50",-- -2827
x"f2b10",-- -3407
x"f1ed0",-- -3603
x"f1090",-- -3831
x"ee470",-- -4537
x"ef3d0",-- -4291
x"f17e0",-- -3714
x"f7ee0",-- -2066
x"fb880",-- -1144
x"fe430",-- -445
x"01380",-- 312
x"03d60",-- 982
x"06d70",-- 1751
x"0ae80",-- 2792
x"0f360",-- 3894
x"12c00",-- 4800
x"14d90",-- 5337
x"167f0",-- 5759
x"18bd0",-- 6333
x"18430",-- 6211
x"198c0",-- 6540
x"1b5a0",-- 7002
x"1c980",-- 7320
x"1c220",-- 7202
x"1b7b0",-- 7035
x"19500",-- 6480
x"19920",-- 6546
x"169a0",-- 5786
x"14750",-- 5237
x"12040",-- 4612
x"146d0",-- 5229
x"17eb0",-- 6123
x"18db0",-- 6363
x"19470",-- 6471
x"18f70",-- 6391
x"1c050",-- 7173
x"1aae0",-- 6830
x"18c00",-- 6336
x"12c20",-- 4802
x"113a0",-- 4410
x"09d10",-- 2513
x"fe110",-- -495
x"eea00",-- -4448
x"e5790",-- -6791
x"e5dd0",-- -6691
x"e9bb0",-- -5701
x"edce0",-- -4658
x"e7d80",-- -6184
x"e05f0",-- -8097
x"dc2d0",-- -9171
x"de710",-- -8591
x"dfc50",-- -8251
x"e3ab0",-- -7253
x"e9d40",-- -5676
x"f0190",-- -4071
x"f5e40",-- -2588
x"fcc60",-- -826
x"01ef0",-- 495
x"02320",-- 562
x"06b80",-- 1720
x"0dc60",-- 3526
x"14a00",-- 5280
x"17a50",-- 6053
x"17cb0",-- 6091
x"14480",-- 5192
x"0e770",-- 3703
x"095d0",-- 2397
x"02580",-- 600
x"fa610",-- -1439
x"f3ba0",-- -3142
x"edb00",-- -4688
x"e5400",-- -6848
x"dd6b0",-- -8853
x"da140",-- -9708
x"d8800",-- -10112
x"d7680",-- -10392
x"d7a90",-- -10327
x"dc0b0",-- -9205
x"e2f00",-- -7440
x"e8710",-- -6031
x"ed650",-- -4763
x"f2060",-- -3578
x"f7f10",-- -2063
x"fd270",-- -729
x"04b80",-- 1208
x"0aa00",-- 2720
x"0d310",-- 3377
x"0e040",-- 3588
x"0f9a0",-- 3994
x"0fdd0",-- 4061
x"0e000",-- 3584
x"0d1c0",-- 3356
x"09fd0",-- 2557
x"05ec0",-- 1516
x"00eb0",-- 235
x"fc3c0",-- -964
x"f5c40",-- -2620
x"f1480",-- -3768
x"ee660",-- -4506
x"eda40",-- -4700
x"ed480",-- -4792
x"edfc0",-- -4612
x"ed5e0",-- -4770
x"ed270",-- -4825
x"f0a50",-- -3931
x"f5dd0",-- -2595
x"fca70",-- -857
x"00b20",-- 178
x"052c0",-- 1324
x"091d0",-- 2333
x"0db70",-- 3511
x"10000",-- 4096
x"11df0",-- 4575
x"13530",-- 4947
x"155f0",-- 5471
x"16fc0",-- 5884
x"18140",-- 6164
x"185c0",-- 6236
x"15ee0",-- 5614
x"15350",-- 5429
x"14860",-- 5254
x"15120",-- 5394
x"154a0",-- 5450
x"14b90",-- 5305
x"131c0",-- 4892
x"12810",-- 4737
x"12270",-- 4647
x"11350",-- 4405
x"0ffb0",-- 4091
x"0fd70",-- 4055
x"12b30",-- 4787
x"166b0",-- 5739
x"1d0f0",-- 7439
x"20b10",-- 8369
x"20320",-- 8242
x"1dab0",-- 7595
x"1b2e0",-- 6958
x"179c0",-- 6044
x"11a50",-- 4517
x"04800",-- 1152
x"f6d90",-- -2343
x"eb0b0",-- -5365
x"e6080",-- -6648
x"e85a0",-- -6054
x"ea290",-- -5591
x"e8260",-- -6106
x"dfc50",-- -8251
x"db7d0",-- -9347
x"dcc40",-- -9020
x"e0370",-- -8137
x"e2760",-- -7562
x"e89e0",-- -5986
x"ee980",-- -4456
x"f5bf0",-- -2625
x"fc710",-- -911
x"02980",-- 664
x"06140",-- 1556
x"08b30",-- 2227
x"0e7c0",-- 3708
x"13790",-- 4985
x"17180",-- 5912
x"17b50",-- 6069
x"15a10",-- 5537
x"10220",-- 4130
x"0a840",-- 2692
x"021c0",-- 540
x"f95e0",-- -1698
x"f12e0",-- -3794
x"eb060",-- -5370
x"e56a0",-- -6806
x"e0330",-- -8141
x"db770",-- -9353
x"d70a0",-- -10486
x"d6870",-- -10617
x"da380",-- -9672
x"e0d50",-- -7979
x"e08f0",-- -8049
x"e1ea0",-- -7702
x"e92a0",-- -5846
x"f78e0",-- -2162
x"03170",-- 791
x"061c0",-- 1564
x"07180",-- 1816
x"09c90",-- 2505
x"0d3d0",-- 3389
x"10cc0",-- 4300
x"13a80",-- 5032
x"0f680",-- 3944
x"0b850",-- 2949
x"08190",-- 2073
x"06d90",-- 1753
x"01b00",-- 432
x"fc0c0",-- -1012
x"f6230",-- -2525
x"f1270",-- -3801
x"edba0",-- -4678
x"eb590",-- -5287
x"e9a10",-- -5727
x"e8ce0",-- -5938
x"ec9d0",-- -4963
x"efce0",-- -4146
x"f3c70",-- -3129
x"f5db0",-- -2597
x"f9700",-- -1680
x"fc620",-- -926
x"02580",-- 600
x"08be0",-- 2238
x"0dc20",-- 3522
x"124d0",-- 4685
x"13380",-- 4920
x"14690",-- 5225
x"14450",-- 5189
x"14b10",-- 5297
x"12f40",-- 4852
x"11860",-- 4486
x"0f8a0",-- 3978
x"0e310",-- 3633
x"0c610",-- 3169
x"0b0e0",-- 2830
x"0a120",-- 2578
x"0a260",-- 2598
x"0bf10",-- 3057
x"0cc80",-- 3272
x"0e3b0",-- 3643
x"0f950",-- 3989
x"11860",-- 4486
x"14930",-- 5267
x"17f80",-- 6136
x"18810",-- 6273
x"18f20",-- 6386
x"1b690",-- 7017
x"22590",-- 8793
x"2a0e0",-- 10766
x"2c510",-- 11345
x"250f0",-- 9487
x"1bdd0",-- 7133
x"15880",-- 5512
x"0dec0",-- 3564
x"ffb50",-- -75
x"f1400",-- -3776
x"e5070",-- -6905
x"dd5f0",-- -8865
x"dcaf0",-- -9041
x"e16b0",-- -7829
x"e1fe0",-- -7682
x"db280",-- -9432
x"d8280",-- -10200
x"dafb0",-- -9477
x"e1860",-- -7802
x"e88a0",-- -6006
x"f1110",-- -3823
x"f7d30",-- -2093
x"ffdb0",-- -37
x"08550",-- 2133
x"0f180",-- 3864
x"12340",-- 4660
x"13f00",-- 5104
x"16be0",-- 5822
x"18e60",-- 6374
x"1a960",-- 6806
x"17c10",-- 6081
x"111a0",-- 4378
x"08c50",-- 2245
x"ffee0",-- -18
x"f5f80",-- -2568
x"ec560",-- -5034
x"e4170",-- -7145
x"dd180",-- -8936
x"d8d00",-- -10032
x"d6ff0",-- -10497
x"d5fc0",-- -10756
x"d5c00",-- -10816
x"d8c90",-- -10039
x"df0a0",-- -8438
x"e7d10",-- -6191
x"f2370",-- -3529
x"fae90",-- -1303
x"01b30",-- 435
x"07010",-- 1793
x"04dc0",-- 1244
x"04340",-- 1076
x"07a30",-- 1955
x"11d20",-- 4562
x"198f0",-- 6543
x"15e70",-- 5607
x"0d5b0",-- 3419
x"03790",-- 889
x"fce60",-- -794
x"fadf0",-- -1313
x"f8410",-- -1983
x"f2b90",-- -3399
x"ef980",-- -4200
x"ea9b0",-- -5477
x"e9bf0",-- -5697
x"e99a0",-- -5734
x"e8460",-- -6074
x"e8e60",-- -5914
x"ead20",-- -5422
x"f1f90",-- -3591
x"f9990",-- -1639
x"ff990",-- -103
x"03f40",-- 1012
x"04d10",-- 1233
x"07ad0",-- 1965
x"0cd20",-- 3282
x"115b0",-- 4443
x"14540",-- 5204
x"14f50",-- 5365
x"134c0",-- 4940
x"11ee0",-- 4590
x"0e070",-- 3591
x"0ae30",-- 2787
x"078d0",-- 1933
x"05b30",-- 1459
x"06520",-- 1618
x"05740",-- 1396
x"056a0",-- 1386
x"03a80",-- 936
x"02780",-- 632
x"04030",-- 1027
x"071f0",-- 1823
x"0bbc0",-- 3004
x"11670",-- 4455
x"17130",-- 5907
x"1dbc0",-- 7612
x"1fd50",-- 8149
x"1f350",-- 7989
x"20450",-- 8261
x"239b0",-- 9115
x"29690",-- 10601
x"2ab50",-- 10933
x"27a30",-- 10147
x"22130",-- 8723
x"1cce0",-- 7374
x"16630",-- 5731
x"09810",-- 2433
x"f4b10",-- -2895
x"e2760",-- -7562
x"d8240",-- -10204
x"d6990",-- -10599
x"da010",-- -9727
x"dcc60",-- -9018
x"dda20",-- -8798
x"db7a0",-- -9350
x"dca60",-- -9050
x"e0e10",-- -7967
x"e7d30",-- -6189
x"f13b0",-- -3781
x"fbd00",-- -1072
x"05260",-- 1318
x"0e8c0",-- 3724
x"15540",-- 5460
x"18660",-- 6246
x"19290",-- 6441
x"18f50",-- 6389
x"189b0",-- 6299
x"176a0",-- 5994
x"15ad0",-- 5549
x"102a0",-- 4138
x"07b30",-- 1971
x"fe410",-- -447
x"f3290",-- -3287
x"e8260",-- -6106
x"df9d0",-- -8291
x"d9500",-- -9904
x"d5b80",-- -10824
x"d5360",-- -10954
x"d6920",-- -10606
x"d8e10",-- -10015
x"dc710",-- -9103
x"e3ab0",-- -7253
x"ec980",-- -4968
x"f7590",-- -2215
x"01810",-- 385
x"099e0",-- 2462
x"0ef40",-- 3828
x"13aa0",-- 5034
x"160f0",-- 5647
x"16bd0",-- 5821
x"159b0",-- 5531
x"09560",-- 2390
x"fead0",-- -339
x"f92a0",-- -1750
x"fe8c0",-- -372
x"014a0",-- 330
x"f9e70",-- -1561
x"ee050",-- -4603
x"e3d30",-- -7213
x"e1b60",-- -7754
x"e5e50",-- -6683
x"e98b0",-- -5749
x"e8cd0",-- -5939
x"eb4d0",-- -5299
x"ed150",-- -4843
x"f5790",-- -2695
x"fc690",-- -919
x"01330",-- 307
x"04ac0",-- 1196
x"072b0",-- 1835
x"0d240",-- 3364
x"11dc0",-- 4572
x"14fa0",-- 5370
x"155d0",-- 5469
x"12d70",-- 4823
x"10040",-- 4100
x"0e0e0",-- 3598
x"09f40",-- 2548
x"074a0",-- 1866
x"01440",-- 324
x"fd3a0",-- -710
x"faeb0",-- -1301
x"fad50",-- -1323
x"fd020",-- -766
x"fda40",-- -604
x"ffcb0",-- -53
x"02780",-- 632
x"05620",-- 1378
x"09e70",-- 2535
x"0e2f0",-- 3631
x"10cf0",-- 4303
x"15080",-- 5384
x"1aa50",-- 6821
x"21600",-- 8544
x"280c0",-- 10252
x"2a520",-- 10834
x"2ad30",-- 10963
x"29f80",-- 10744
x"28b60",-- 10422
x"27e40",-- 10212
x"1fc30",-- 8131
x"17710",-- 6001
x"12140",-- 4628
x"0b530",-- 2899
x"fbf60",-- -1034
x"e9660",-- -5786
x"d8f00",-- -10000
x"cff50",-- -12299
x"ceba0",-- -12614
x"d8130",-- -10221
x"e1fc0",-- -7684
x"e3c90",-- -7223
x"e4b40",-- -6988
x"e7e70",-- -6169
x"ee800",-- -4480
x"f5c50",-- -2619
x"feca0",-- -310
x"07090",-- 1801
x"0ed10",-- 3793
x"17b50",-- 6069
x"1d8c0",-- 7564
x"1cdb0",-- 7387
x"19120",-- 6418
x"14570",-- 5207
x"0eed0",-- 3821
x"0ceb0",-- 3307
x"0a400",-- 2624
x"04670",-- 1127
x"fb5b0",-- -1189
x"f2170",-- -3561
x"e8230",-- -6109
x"de080",-- -8696
x"d8a50",-- -10075
x"d5f50",-- -10763
x"d6920",-- -10606
x"db320",-- -9422
x"e10a0",-- -7926
x"e6780",-- -6536
x"ec6c0",-- -5012
x"f2f50",-- -3339
x"faf00",-- -1296
x"04390",-- 1081
x"0dfa0",-- 3578
x"14340",-- 5172
x"17560",-- 5974
x"180f0",-- 6159
x"14f90",-- 5369
x"10590",-- 4185
x"0c080",-- 3080
x"05f30",-- 1523
x"ff560",-- -170
x"f7750",-- -2187
x"e75c0",-- -6308
x"db900",-- -9328
x"dcf50",-- -8971
x"e7840",-- -6268
x"ecad0",-- -4947
x"e9d90",-- -5671
x"e7c20",-- -6206
x"e94d0",-- -5811
x"ee1a0",-- -4582
x"f6370",-- -2505
x"fbb70",-- -1097
x"fe2b0",-- -469
x"042b0",-- 1067
x"0b440",-- 2884
x"12a70",-- 4775
x"16980",-- 5784
x"14ed0",-- 5357
x"0ed40",-- 3796
x"0afc0",-- 2812
x"0b170",-- 2839
x"0c180",-- 3096
x"0ae50",-- 2789
x"07680",-- 1896
x"01db0",-- 475
x"fc8e0",-- -882
x"f9830",-- -1661
x"f4120",-- -3054
x"f1c90",-- -3639
x"f3b60",-- -3146
x"faf00",-- -1296
x"00780",-- 120
x"03ae0",-- 942
x"05420",-- 1346
x"072c0",-- 1836
x"0b600",-- 2912
x"13360",-- 4918
x"19350",-- 6453
x"1d230",-- 7459
x"1f960",-- 8086
x"216e0",-- 8558
x"26bb0",-- 9915
x"2afc0",-- 11004
x"2d7f0",-- 11647
x"2a720",-- 10866
x"26ba0",-- 9914
x"24200",-- 9248
x"1dda0",-- 7642
x"11df0",-- 4575
x"06000",-- 1536
x"fa140",-- -1516
x"ed9d0",-- -4707
x"dd610",-- -8863
x"cf450",-- -12475
x"cc740",-- -13196
x"d4d80",-- -11048
x"e2f60",-- -7434
x"e9bb0",-- -5701
x"e88a0",-- -6006
x"e8830",-- -6013
x"ef6d0",-- -4243
x"f8ff0",-- -1793
x"02a70",-- 679
x"0a2d0",-- 2605
x"10810",-- 4225
x"15540",-- 5460
x"1ad10",-- 6865
x"1db50",-- 7605
x"1a8e0",-- 6798
x"14e00",-- 5344
x"0e2d0",-- 3629
x"095d0",-- 2397
x"06c70",-- 1735
x"03c90",-- 969
x"fc2a0",-- -982
x"f1fe0",-- -3586
x"e8850",-- -6011
x"e0d80",-- -7976
x"daf10",-- -9487
x"d8c10",-- -10047
x"d9360",-- -9930
x"dbf60",-- -9226
x"e30a0",-- -7414
x"eac60",-- -5434
x"f1cf0",-- -3633
x"f8d50",-- -1835
x"00210",-- 33
x"073b0",-- 1851
x"0e680",-- 3688
x"14e00",-- 5344
x"17af0",-- 6063
x"16fa0",-- 5882
x"14410",-- 5185
x"0eff0",-- 3839
x"092c0",-- 2348
x"02e00",-- 736
x"fc340",-- -972
x"f5340",-- -2764
x"ef770",-- -4233
x"ebcc0",-- -5172
x"e77c0",-- -6276
x"e6500",-- -6576
x"e1e20",-- -7710
x"de010",-- -8703
x"daeb0",-- -9493
x"e2550",-- -7595
x"ef600",-- -4256
x"fb4f0",-- -1201
x"02ed0",-- 749
x"04340",-- 1076
x"06690",-- 1641
x"09580",-- 2392
x"0e1e0",-- 3614
x"116f0",-- 4463
x"13260",-- 4902
x"11c30",-- 4547
x"11330",-- 4403
x"0f580",-- 3928
x"0c9f0",-- 3231
x"072b0",-- 1835
x"005d0",-- 93
x"fb3b0",-- -1221
x"f8440",-- -1980
x"f8960",-- -1898
x"f9070",-- -1785
x"f8230",-- -2013
x"f7330",-- -2253
x"f8390",-- -1991
x"fa390",-- -1479
x"feed0",-- -275
x"033a0",-- 826
x"07f10",-- 2033
x"0b3a0",-- 2874
x"0d1a0",-- 3354
x"0ffa0",-- 4090
x"13fb0",-- 5115
x"19830",-- 6531
x"1d460",-- 7494
x"1f1c0",-- 7964
x"203c0",-- 8252
x"218d0",-- 8589
x"229c0",-- 8860
x"21d30",-- 8659
x"20390",-- 8249
x"205c0",-- 8284
x"21ba0",-- 8634
x"1fb20",-- 8114
x"1a910",-- 6801
x"0bee0",-- 3054
x"ef700",-- -4240
x"cf960",-- -12394
x"c2180",-- -15848
x"cd2f0",-- -13009
x"df540",-- -8364
x"ec6c0",-- -5012
x"efa40",-- -4188
x"ef610",-- -4255
x"eec60",-- -4410
x"f2df0",-- -3361
x"f5770",-- -2697
x"f7fd0",-- -2051
x"fe850",-- -379
x"0a8e0",-- 2702
x"18110",-- 6161
x"21740",-- 8564
x"220a0",-- 8714
x"184d0",-- 6221
x"0d1c0",-- 3356
x"065f0",-- 1631
x"05c70",-- 1479
x"073b0",-- 1851
x"07ea0",-- 2026
x"03a40",-- 932
x"fb5e0",-- -1186
x"f1450",-- -3771
x"e5e20",-- -6686
x"db430",-- -9405
x"d5610",-- -10911
x"d6c60",-- -10554
x"dde30",-- -8733
x"e7ca0",-- -6198
x"efd90",-- -4135
x"f4620",-- -2974
x"f7db0",-- -2085
x"fca20",-- -862
x"03040",-- 772
x"0aeb0",-- 2795
x"12d60",-- 4822
x"178c0",-- 6028
x"18d20",-- 6354
x"167f0",-- 5759
x"10870",-- 4231
x"07e90",-- 2025
x"fef70",-- -265
x"f7fd0",-- -2051
x"f28c0",-- -3444
x"f09e0",-- -3938
x"ef420",-- -4286
x"edb80",-- -4680
x"ea920",-- -5486
x"e82d0",-- -6099
x"e6c10",-- -6463
x"e9cf0",-- -5681
x"ec8f0",-- -4977
x"ea3d0",-- -5571
x"ecdf0",-- -4897
x"f2100",-- -3568
x"fe2b0",-- -469
x"08630",-- 2147
x"0e1d0",-- 3613
x"0fe20",-- 4066
x"0cc80",-- 3272
x"0d400",-- 3392
x"0f8f0",-- 3983
x"0f120",-- 3858
x"0deb0",-- 3563
x"0aca0",-- 2762
x"05720",-- 1394
x"03920",-- 914
x"011f0",-- 287
x"fdf10",-- -527
x"f9090",-- -1783
x"f3950",-- -3179
x"f2ac0",-- -3412
x"f44d0",-- -2995
x"f8610",-- -1951
x"fcc80",-- -824
x"fe0c0",-- -500
x"008a0",-- 138
x"03810",-- 897
x"06b30",-- 1715
x"0b220",-- 2850
x"0e500",-- 3664
x"10d70",-- 4311
x"12960",-- 4758
x"13c90",-- 5065
x"14200",-- 5152
x"10de0",-- 4318
x"10590",-- 4185
x"12430",-- 4675
x"17e60",-- 6118
x"1c4a0",-- 7242
x"1db20",-- 7602
x"1c930",-- 7315
x"1aa70",-- 6823
x"196e0",-- 6510
x"1b100",-- 6928
x"1d910",-- 7569
x"1be90",-- 7145
x"0cc30",-- 3267
x"e9680",-- -5784
x"ca9a0",-- -13670
x"c6300",-- -14800
x"dbc20",-- -9278
x"ee5d0",-- -4515
x"f3610",-- -3231
x"f1c40",-- -3644
x"f0a50",-- -3931
x"f2390",-- -3527
x"f5650",-- -2715
x"f6200",-- -2528
x"f49b0",-- -2917
x"f8d00",-- -1840
x"059e0",-- 1438
x"164f0",-- 5711
x"21d00",-- 8656
x"22600",-- 8800
x"167a0",-- 5754
x"09900",-- 2448
x"03e70",-- 999
x"050e0",-- 1294
x"07e00",-- 2016
x"08170",-- 2071
x"03620",-- 866
x"fb090",-- -1271
x"f19d0",-- -3683
x"e6960",-- -6506
x"dabc0",-- -9540
x"d4a80",-- -11096
x"d7770",-- -10377
x"e0290",-- -8151
x"eae30",-- -5405
x"f4550",-- -2987
x"fa110",-- -1519
x"fd1f0",-- -737
x"00be0",-- 190
x"04dc0",-- 1244
x"0b0e0",-- 2830
x"11bf0",-- 4543
x"16230",-- 5667
x"16c50",-- 5829
x"14d70",-- 5335
x"0f8d0",-- 3981
x"06bb0",-- 1723
x"fd760",-- -650
x"f5a70",-- -2649
x"f1390",-- -3783
x"efdb0",-- -4133
x"f0710",-- -3983
x"ef450",-- -4283
x"ecaf0",-- -4945
x"ea620",-- -5534
x"e88d0",-- -6003
x"e98e0",-- -5746
x"ee010",-- -4607
x"f5570",-- -2729
x"fcc00",-- -832
x"05310",-- 1329
x"08580",-- 2136
x"07760",-- 1910
x"05e70",-- 1511
x"05a90",-- 1449
x"034a0",-- 842
x"02670",-- 615
x"06e00",-- 1760
x"0d240",-- 3364
x"0f8d0",-- 3981
x"0b9a0",-- 2970
x"05790",-- 1401
x"fdc20",-- -574
x"f9330",-- -1741
x"f76a0",-- -2198
x"f7770",-- -2185
x"f8850",-- -1915
x"fadc0",-- -1316
x"fbdd0",-- -1059
x"fd2e0",-- -722
x"fd0b0",-- -757
x"fcc80",-- -824
x"fd800",-- -640
x"ff800",-- -128
x"04d90",-- 1241
x"0a000",-- 2560
x"0de70",-- 3559
x"0f060",-- 3846
x"0d630",-- 3427
x"0c430",-- 3139
x"0b800",-- 2944
x"0a5f0",-- 2655
x"07ab0",-- 1963
x"042a0",-- 1066
x"03760",-- 886
x"06730",-- 1651
x"0b810",-- 2945
x"0da80",-- 3496
x"0e2c0",-- 3628
x"0d270",-- 3367
x"0f6d0",-- 3949
x"11dc0",-- 4572
x"17b00",-- 6064
x"1cf40",-- 7412
x"24470",-- 9287
x"28ab0",-- 10411
x"2d620",-- 11618
x"29490",-- 10569
x"f6190",-- -2535
x"c1840",-- -15996
x"b5160",-- -19178
x"d6ff0",-- -10497
x"ef980",-- -4200
x"f3810",-- -3199
x"f4940",-- -2924
x"f0c80",-- -3896
x"ef340",-- -4300
x"f4730",-- -2957
x"f5bf0",-- -2625
x"ef5e0",-- -4258
x"f21e0",-- -3554
x"00700",-- 112
x"17290",-- 5929
x"2b2b0",-- 11051
x"31f70",-- 12791
x"1f120",-- 7954
x"06f70",-- 1783
x"faeb0",-- -1301
x"f9c90",-- -1591
x"fdcb0",-- -565
x"02890",-- 649
x"01170",-- 279
x"fc440",-- -956
x"f7b50",-- -2123
x"ee0d0",-- -4595
x"ddf60",-- -8714
x"d35e0",-- -11426
x"d5020",-- -11006
x"dc870",-- -9081
x"eafc0",-- -5380
x"fb360",-- -1226
x"047b0",-- 1147
x"06b30",-- 1715
x"05920",-- 1426
x"04cd0",-- 1229
x"07130",-- 1811
x"0d400",-- 3392
x"119a0",-- 4506
x"13870",-- 4999
x"15fd0",-- 5629
x"146d0",-- 5229
x"0b6c0",-- 2924
x"ffe50",-- -27
x"f4280",-- -3032
x"ea830",-- -5501
x"e7340",-- -6348
x"e8e10",-- -5919
x"ea650",-- -5531
x"ea650",-- -5531
x"eb470",-- -5305
x"eb110",-- -5359
x"ed390",-- -4807
x"f3040",-- -3324
x"fa170",-- -1513
x"01630",-- 355
x"0a0a0",-- 2570
x"11df0",-- 4575
x"16f00",-- 5872
x"19350",-- 6453
x"17220",-- 5922
x"13590",-- 4953
x"0d1c0",-- 3356
x"021c0",-- 540
x"f72c0",-- -2260
x"f5f40",-- -2572
x"f9ae0",-- -1618
x"f9bf0",-- -1601
x"f7da0",-- -2086
x"f71a0",-- -2278
x"f7630",-- -2205
x"f6120",-- -2542
x"f66b0",-- -2453
x"f6a20",-- -2398
x"f74f0",-- -2225
x"fb420",-- -1214
x"ff3a0",-- -198
x"03bf0",-- 959
x"08a00",-- 2208
x"09510",-- 2385
x"08480",-- 2120
x"06d60",-- 1750
x"06ea0",-- 1770
x"06700",-- 1648
x"061b0",-- 1563
x"065a0",-- 1626
x"060c0",-- 1548
x"05bc0",-- 1468
x"04fe0",-- 1278
x"01ef0",-- 495
x"fea20",-- -350
x"fdfd0",-- -515
x"fecb0",-- -309
x"00e80",-- 232
x"02800",-- 640
x"035e0",-- 862
x"03310",-- 817
x"04c20",-- 1218
x"069b0",-- 1691
x"08870",-- 2183
x"0ae10",-- 2785
x"0cd20",-- 3282
x"108e0",-- 4238
x"14480",-- 5192
x"19bf0",-- 6591
x"1d3d0",-- 7485
x"1fc60",-- 8134
x"1fdf0",-- 8159
x"20f40",-- 8436
x"20160",-- 8214
x"0c7d0",-- 3197
x"e9480",-- -5816
x"cbe10",-- -13343
x"cc4e0",-- -13234
x"dcd00",-- -9008
x"ed1a0",-- -4838
x"f4370",-- -3017
x"f4fd0",-- -2819
x"f40d0",-- -3059
x"f6080",-- -2552
x"f81c0",-- -2020
x"f6af0",-- -2385
x"f4dc0",-- -2852
x"f6200",-- -2528
x"ff1c0",-- -228
x"0e570",-- 3671
x"1ce50",-- 7397
x"1e4d0",-- 7757
x"13310",-- 4913
x"05950",-- 1429
x"fd850",-- -635
x"fd450",-- -699
x"00760",-- 118
x"02fc0",-- 764
x"02550",-- 597
x"008a0",-- 138
x"fc0d0",-- -1011
x"f3180",-- -3304
x"e8e40",-- -5916
x"e0990",-- -8039
x"ddbd0",-- -8771
x"e1970",-- -7785
x"eb4f0",-- -5297
x"f6760",-- -2442
x"ff1f0",-- -225
x"034c0",-- 844
x"03f10",-- 1009
x"049b0",-- 1179
x"07a90",-- 1961
x"0b3a0",-- 2874
x"0e020",-- 3586
x"0fff0",-- 4095
x"0f310",-- 3889
x"0ade0",-- 2782
x"04840",-- 1156
x"fce40",-- -796
x"f4e60",-- -2842
x"ee700",-- -4496
x"ebd80",-- -5160
x"ebcf0",-- -5169
x"ee980",-- -4456
x"f2010",-- -3583
x"f4c00",-- -2880
x"f6d70",-- -2345
x"f9970",-- -1641
x"fd670",-- -665
x"020a0",-- 522
x"07e40",-- 2020
x"0cdc0",-- 3292
x"103e0",-- 4158
x"131a0",-- 4890
x"13bc0",-- 5052
x"11d50",-- 4565
x"0dd30",-- 3539
x"09bf0",-- 2495
x"05950",-- 1429
x"02570",-- 599
x"000f0",-- 15
x"fe5d0",-- -419
x"f8490",-- -1975
x"ef1a0",-- -4326
x"e96b0",-- -5781
x"eb0c0",-- -5364
x"f0260",-- -4058
x"f0760",-- -3978
x"f1fb0",-- -3589
x"f5ef0",-- -2577
x"fc300",-- -976
x"00c50",-- 197
x"02af0",-- 687
x"03e40",-- 996
x"05830",-- 1411
x"086e0",-- 2158
x"0c6b0",-- 3179
x"0f130",-- 3859
x"0f7b0",-- 3963
x"0b770",-- 2935
x"05220",-- 1314
x"008f0",-- 143
x"fdfe0",-- -514
x"fb4f0",-- -1201
x"f9070",-- -1785
x"f8be0",-- -1858
x"fa0a0",-- -1526
x"fc110",-- -1007
x"fc690",-- -919
x"fb850",-- -1147
x"faca0",-- -1334
x"fc780",-- -904
x"fffd0",-- -3
x"03bd0",-- 957
x"08820",-- 2178
x"0c9b0",-- 3227
x"0ea20",-- 3746
x"0f040",-- 3844
x"0eae0",-- 3758
x"0e9a0",-- 3738
x"0f300",-- 3888
x"104f0",-- 4175
x"12e80",-- 4840
x"151a0",-- 5402
x"17bc0",-- 6076
x"16ca0",-- 5834
x"16630",-- 5731
x"15850",-- 5509
x"14ed0",-- 5357
x"0c180",-- 3096
x"f5ca0",-- -2614
x"dc460",-- -9146
x"d0150",-- -12267
x"d9730",-- -9869
x"e8350",-- -6091
x"f33e0",-- -3266
x"f7360",-- -2250
x"f90b0",-- -1781
x"f9990",-- -1639
x"fa710",-- -1423
x"fa910",-- -1391
x"f9100",-- -1776
x"f7b80",-- -2120
x"fbd60",-- -1066
x"06250",-- 1573
x"15210",-- 5409
x"1e1d0",-- 7709
x"1b7b0",-- 7035
x"10520",-- 4178
x"05df0",-- 1503
x"00870",-- 135
x"feeb0",-- -277
x"fedf0",-- -289
x"febb0",-- -325
x"fd950",-- -619
x"fb8d0",-- -1139
x"f6d70",-- -2345
x"ef920",-- -4206
x"e8300",-- -6096
x"e1ac0",-- -7764
x"e05b0",-- -8101
x"e5e80",-- -6680
x"f19f0",-- -3681
x"fdea0",-- -534
x"06610",-- 1633
x"0a640",-- 2660
x"0a860",-- 2694
x"08320",-- 2098
x"05c70",-- 1479
x"058b0",-- 1419
x"06a50",-- 1701
x"091d0",-- 2333
x"0b5d0",-- 2909
x"0b600",-- 2912
x"085e0",-- 2142
x"01bd0",-- 445
x"f9b30",-- -1613
x"f2780",-- -3464
x"efb80",-- -4168
x"f10c0",-- -3828
x"f4f80",-- -2824
x"f8ee0",-- -1810
x"fc030",-- -1021
x"fd670",-- -665
x"fdd10",-- -559
x"fd9c0",-- -612
x"fdfd0",-- -515
x"fff30",-- -13
x"03d60",-- 982
x"08c50",-- 2245
x"0d590",-- 3417
x"0fdd0",-- 4061
x"0f450",-- 3909
x"0bf10",-- 3057
x"078a0",-- 1930
x"03ba0",-- 954
x"01490",-- 329
x"00670",-- 103
x"001c0",-- 28
x"ff950",-- -107
x"fe780",-- -392
x"fccb0",-- -821
x"fa6b0",-- -1429
x"f8070",-- -2041
x"f6730",-- -2445
x"f6750",-- -2443
x"f8bb0",-- -1861
x"fc170",-- -1001
x"ffcb0",-- -53
x"02b10",-- 689
x"04fa0",-- 1274
x"05fd0",-- 1533
x"06d20",-- 1746
x"07630",-- 1891
x"07d00",-- 2000
x"08030",-- 2051
x"07cc0",-- 1996
x"06f20",-- 1778
x"05120",-- 1298
x"02210",-- 545
x"fe7b0",-- -389
x"faaf0",-- -1361
x"f7ee0",-- -2066
x"f4bc0",-- -2884
x"efa40",-- -4188
x"ed1f0",-- -4833
x"ed510",-- -4783
x"edd60",-- -4650
x"edd90",-- -4647
x"f0d00",-- -3888
x"f6b10",-- -2383
x"fb9e0",-- -1122
x"fe460",-- -442
x"00870",-- 135
x"01030",-- 259
x"02480",-- 584
x"03e50",-- 997
x"04dc0",-- 1244
x"064d0",-- 1613
x"06b10",-- 1713
x"064e0",-- 1614
x"04a50",-- 1189
x"030e0",-- 782
x"01790",-- 377
x"fdf40",-- -524
x"faf50",-- -1291
x"f9fb0",-- -1541
x"fb6d0",-- -1171
x"feac0",-- -340
x"01f80",-- 504
x"047d0",-- 1149
x"05e20",-- 1506
x"07380",-- 1848
x"07860",-- 1926
x"08500",-- 2128
x"093b0",-- 2363
x"0b830",-- 2947
x"0e570",-- 3671
x"14220",-- 5154
x"1a750",-- 6773
x"21210",-- 8481
x"24bd0",-- 9405
x"29320",-- 10546
x"2f580",-- 12120
x"300b0",-- 12299
x"1a5e0",-- 6750
x"e5b30",-- -6733
x"c4330",-- -15309
x"c60e0",-- -14834
x"dd720",-- -8846
x"e95e0",-- -5794
x"ec710",-- -5007
x"f1c20",-- -3646
x"f40d0",-- -3059
x"f9700",-- -1680
x"fb400",-- -1216
x"f6b40",-- -2380
x"ef4d0",-- -4275
x"eb5b0",-- -5285
x"f6730",-- -2445
x"10780",-- 4216
x"2d960",-- 11670
x"36c90",-- 14025
x"27920",-- 10130
x"149f0",-- 5279
x"07400",-- 1856
x"024e0",-- 590
x"fe390",-- -455
x"fc750",-- -907
x"fc030",-- -1021
x"fd400",-- -704
x"005d0",-- 93
x"fe500",-- -432
x"f5790",-- -2695
x"e7520",-- -6318
x"d7390",-- -10439
x"d1140",-- -12012
x"d90c0",-- -9972
x"ec350",-- -5067
x"fd720",-- -654
x"085c0",-- 2140
x"0de50",-- 3557
x"10550",-- 4181
x"11580",-- 4440
x"0ebe0",-- 3774
x"0b240",-- 2852
x"08f00",-- 2288
x"0a390",-- 2617
x"0f310",-- 3889
x"13ec0",-- 5100
x"14360",-- 5174
x"0b880",-- 2952
x"fcb60",-- -842
x"eedc0",-- -4388
x"e6ff0",-- -6401
x"e5a70",-- -6745
x"e6af0",-- -6481
x"e96a0",-- -5782
x"ee3c0",-- -4548
x"f3f30",-- -3085
x"f96d0",-- -1683
x"fd1d0",-- -739
x"fdb00",-- -592
x"fcf30",-- -781
x"fe700",-- -400
x"04700",-- 1136
x"0cd90",-- 3289
x"14e30",-- 5347
x"18b80",-- 6328
x"173c0",-- 5948
x"132c0",-- 4908
x"0e370",-- 3639
x"08a70",-- 2215
x"029e0",-- 670
x"fcda0",-- -806
x"f8520",-- -1966
x"f6550",-- -2475
x"f70c0",-- -2292
x"f76f0",-- -2193
x"f5010",-- -2815
x"f12f0",-- -3793
x"edb30",-- -4685
x"edf90",-- -4615
x"f20a0",-- -3574
x"f8260",-- -2010
x"fdf60",-- -522
x"02e00",-- 736
x"08930",-- 2195
x"0cbd0",-- 3261
x"0ff60",-- 4086
x"10250",-- 4133
x"0e0f0",-- 3599
x"0b260",-- 2854
x"08ca0",-- 2250
x"079c0",-- 1948
x"05fb0",-- 1531
x"031d0",-- 797
x"febb0",-- -325
x"fa000",-- -1536
x"f6580",-- -2472
x"f3390",-- -3271
x"f0c50",-- -3899
x"ef380",-- -4296
x"eeb10",-- -4431
x"f0800",-- -3968
x"f4250",-- -3035
x"f9010",-- -1791
x"fd4a0",-- -694
x"00b60",-- 182
x"03630",-- 867
x"061b0",-- 1563
x"095e0",-- 2398
x"0ba40",-- 2980
x"0c950",-- 3221
x"0cbb0",-- 3259
x"0be20",-- 3042
x"0a9a0",-- 2714
x"08170",-- 2071
x"04b30",-- 1203
x"003f0",-- 63
x"fb8a0",-- -1142
x"f7ce0",-- -2098
x"f5560",-- -2730
x"f4aa0",-- -2902
x"f4d50",-- -2859
x"f5310",-- -2767
x"f7360",-- -2250
x"f9ba0",-- -1606
x"fbf90",-- -1031
x"fdba0",-- -582
x"ff220",-- -222
x"00570",-- 87
x"017b0",-- 379
x"03fe0",-- 1022
x"06860",-- 1670
x"087d0",-- 2173
x"09920",-- 2450
x"09900",-- 2448
x"09180",-- 2328
x"078a0",-- 1930
x"055d0",-- 1373
x"02ca0",-- 714
x"007d0",-- 125
x"feb20",-- -334
x"fd070",-- -761
x"fca20",-- -862
x"fc4d0",-- -947
x"fb520",-- -1198
x"fa1c0",-- -1508
x"f8fc0",-- -1796
x"f8f70",-- -1801
x"f9c20",-- -1598
x"fbd30",-- -1069
x"fe490",-- -439
x"01620",-- 354
x"04d40",-- 1236
x"07710",-- 1905
x"08a70",-- 2215
x"07ef0",-- 2031
x"045a0",-- 1114
x"002f0",-- 47
x"fdc90",-- -567
x"fde90",-- -535
x"ff600",-- -160
x"00af0",-- 175
x"01380",-- 312
x"00bc0",-- 188
x"00050",-- 5
x"ff3d0",-- -195
x"fe530",-- -429
x"fd880",-- -632
x"fd600",-- -672
x"fe210",-- -479
x"007d0",-- 125
x"02c10",-- 705
x"03ba0",-- 954
x"02690",-- 617
x"00940",-- 148
x"fef30",-- -269
x"febb0",-- -325
x"ffdf0",-- -33
x"01770",-- 375
x"03120",-- 786
x"03fb0",-- 1019
x"04d40",-- 1236
x"04b10",-- 1201
x"03a30",-- 931
x"01710",-- 369
x"ff260",-- -218
x"fde00",-- -544
x"fe1b0",-- -485
x"ff510",-- -175
x"ffe70",-- -25
x"ff950",-- -107
x"fe870",-- -377
x"fd710",-- -655
x"fcbb0",-- -837
x"fc700",-- -912
x"fc850",-- -891
x"fcd00",-- -816
x"fde40",-- -540
x"ffa40",-- -92
x"01290",-- 297
x"020f0",-- 527
x"02260",-- 550
x"01df0",-- 479
x"01380",-- 312
x"01790",-- 377
x"fe5d0",-- -419
x"f92a0",-- -1750
x"f5880",-- -2680
x"f5a90",-- -2647
x"f8de0",-- -1826
x"fa930",-- -1389
x"fc6b0",-- -917
x"fc000",-- -1024
x"fb2a0",-- -1238
x"f9f60",-- -1546
x"f8160",-- -2026
x"f8370",-- -1993
x"f8aa0",-- -1878
x"f92a0",-- -1750
x"fa850",-- -1403
x"fe020",-- -510
x"03620",-- 866
x"05f60",-- 1526
x"067d0",-- 1661
x"05770",-- 1399
x"04710",-- 1137
x"05090",-- 1289
x"06350",-- 1589
x"093a0",-- 2362
x"0e3e0",-- 3646
x"132e0",-- 4910
x"163c0",-- 5692
x"169b0",-- 5787
x"16960",-- 5782
x"15910",-- 5521
x"14090",-- 5129
x"13760",-- 4982
x"13440",-- 4932
x"117e0",-- 4478
x"07c70",-- 1991
x"f71a0",-- -2278
x"e91f0",-- -5857
x"e59d0",-- -6755
x"e7fc0",-- -6148
x"e9ef0",-- -5649
x"ebbd0",-- -5187
x"ef3e0",-- -4290
x"f34a0",-- -3254
x"f76f0",-- -2193
x"fa1e0",-- -1506
x"fa200",-- -1504
x"f7740",-- -2188
x"f3f40",-- -3084
x"f3a60",-- -3162
x"faff0",-- -1281
x"08160",-- 2070
x"12d90",-- 4825
x"17730",-- 6003
x"17a30",-- 6051
x"159b0",-- 5531
x"12780",-- 4728
x"0e980",-- 3736
x"09e00",-- 2528
x"04dc0",-- 1244
x"00070",-- 7
x"fca70",-- -857
x"faf20",-- -1294
x"fac50",-- -1339
x"f90e0",-- -1778
x"f3610",-- -3231
x"eb9c0",-- -5220
x"e57a0",-- -6790
x"e3db0",-- -7205
x"e6730",-- -6541
x"eb790",-- -5255
x"f16b0",-- -3733
x"f7560",-- -2218
x"fd8a0",-- -630
x"03030",-- 771
x"080f0",-- 2063
x"0bab0",-- 2987
x"0c5e0",-- 3166
x"0abb0",-- 2747
x"09210",-- 2337
x"09b00",-- 2480
x"0b720",-- 2930
x"0cbd0",-- 3261
x"0c310",-- 3121
x"097c0",-- 2428
x"056f0",-- 1391
x"00af0",-- 175
x"fbec0",-- -1044
x"f7430",-- -2237
x"f2f70",-- -3337
x"ef750",-- -4235
x"ede30",-- -4637
x"ef4d0",-- -4275
x"f2e80",-- -3352
x"f6bc0",-- -2372
x"f94c0",-- -1716
x"fa780",-- -1416
x"fb880",-- -1144
x"fd770",-- -649
x"00170",-- 23
x"02fa0",-- 762
x"05d10",-- 1489
x"08a50",-- 2213
x"0b1d0",-- 2845
x"0d290",-- 3369
x"0e610",-- 3681
x"0e4b0",-- 3659
x"0cbd0",-- 3261
x"09650",-- 2405
x"05830",-- 1411
x"02410",-- 577
x"00490",-- 73
x"ff4a0",-- -182
x"fe5d0",-- -419
x"fd470",-- -697
x"fbe40",-- -1052
x"fa8f0",-- -1393
x"f9a10",-- -1631
x"f8fd0",-- -1795
x"f8550",-- -1963
x"f7950",-- -2155
x"f74f0",-- -2225
x"f84e0",-- -1970
x"fa9d0",-- -1379
x"fda40",-- -604
x"fffb0",-- -5
x"014e0",-- 334
x"02200",-- 544
x"03210",-- 801
x"042d0",-- 1069
x"051a0",-- 1306
x"05950",-- 1429
x"05510",-- 1361
x"04b80",-- 1208
x"04500",-- 1104
x"047a0",-- 1146
x"04980",-- 1176
x"04490",-- 1097
x"02eb0",-- 747
x"00f90",-- 249
x"ff180",-- -232
x"fd8b0",-- -629
x"fc2d0",-- -979
x"fafa0",-- -1286
x"f9d80",-- -1576
x"f9110",-- -1775
x"f91a0",-- -1766
x"f9bf0",-- -1601
x"faa70",-- -1369
x"fb670",-- -1177
x"fc1c0",-- -996
x"fca80",-- -856
x"fd720",-- -654
x"feb90",-- -327
x"001b0",-- 27
x"018a0",-- 394
x"030e0",-- 782
x"048a0",-- 1162
x"05ef0",-- 1519
x"06c30",-- 1731
x"06d20",-- 1746
x"05e90",-- 1513
x"04b60",-- 1206
x"03490",-- 841
x"02000",-- 512
x"01310",-- 305
x"00c10",-- 193
x"00610",-- 97
x"00000",-- 0
x"ff900",-- -112
x"feed0",-- -275
x"fe1b0",-- -485
x"fd100",-- -752
x"fc0a0",-- -1014
x"fb3e0",-- -1218
x"fb400",-- -1216
x"fbee0",-- -1042
x"fd1a0",-- -742
x"fe690",-- -407
x"ffb20",-- -78
x"00a00",-- 160
x"01990",-- 409
x"02670",-- 615
x"02fa0",-- 762
x"03670",-- 871
x"03d30",-- 979
x"04410",-- 1089
x"04a50",-- 1189
x"04910",-- 1169
x"03620",-- 866
x"016d0",-- 365
x"ffc40",-- -60
x"feb10",-- -335
x"fe3a0",-- -454
x"fe120",-- -494
x"fe140",-- -492
x"fe580",-- -424
x"feeb0",-- -277
x"ffd10",-- -47
x"00820",-- 130
x"00eb0",-- 235
x"00c50",-- 197
x"00580",-- 88
x"00610",-- 97
x"00cf0",-- 207
x"01350",-- 309
x"01270",-- 295
x"00eb0",-- 235
x"00a00",-- 160
x"00370",-- 55
x"00500",-- 80
x"008c0",-- 140
x"00b20",-- 178
x"00cf0",-- 207
x"00fc0",-- 252
x"016d0",-- 365
x"01fb0",-- 507
x"025c0",-- 604
x"023e0",-- 574
x"01db0",-- 475
x"01a30",-- 419
x"01760",-- 374
x"016a0",-- 362
x"01620",-- 354
x"01290",-- 297
x"00f40",-- 244
x"00b60",-- 182
x"00aa0",-- 170
x"00930",-- 147
x"005f0",-- 95
x"000f0",-- 15
x"ffbf0",-- -65
x"ff880",-- -120
x"ff850",-- -123
x"ffc60",-- -58
x"00210",-- 33
x"00390",-- 57
x"00160",-- 22
x"ffe00",-- -32
x"ffa30",-- -93
x"ff6c0",-- -148
x"ff290",-- -215
x"ff0c0",-- -244
x"ff040",-- -252
x"ff0c0",-- -244
x"ff150",-- -235
x"ff3b0",-- -197
x"ff950",-- -107
x"00000",-- 0
x"00800",-- 128
x"00fe0",-- 254
x"01810",-- 385
x"01df0",-- 479
x"02350",-- 565
x"025c0",-- 604
x"025f0",-- 607
x"023c0",-- 572
x"021e0",-- 542
x"01d00",-- 464
x"014c0",-- 332
x"00d50",-- 213
x"00480",-- 72
x"ff8d0",-- -115
x"fe930",-- -365
x"fdc90",-- -567
x"fd3a0",-- -710
x"fcfc0",-- -772
x"fcd40",-- -812
x"fced0",-- -787
x"fd3d0",-- -707
x"fd990",-- -615
x"fe0f0",-- -497
x"fe8f0",-- -369
x"ff070",-- -249
x"ff7c0",-- -132
x"fffb0",-- -5
x"00960",-- 150
x"017b0",-- 379
x"023c0",-- 572
x"029d0",-- 669
x"02af0",-- 687
x"029b0",-- 667
x"02610",-- 609
x"02120",-- 530
x"01a30",-- 419
x"01180",-- 280
x"009e0",-- 158
x"00250",-- 37
x"ffa60",-- -90
x"ff0b0",-- -245
x"fe8e0",-- -370
x"fe140",-- -492
x"fdb30",-- -589
x"fdb20",-- -590
x"fdda0",-- -550
x"fe430",-- -445
x"fea50",-- -347
x"fed40",-- -300
x"fefa0",-- -262
x"fefd0",-- -259
x"ff060",-- -250
x"ff040",-- -252
x"ff310",-- -207
x"ffab0",-- -85
x"00140",-- 20
x"007a0",-- 122
x"00c50",-- 197
x"00fc0",-- 252
x"01150",-- 277
x"01040",-- 260
x"00f50",-- 245
x"00eb0",-- 235
x"01150",-- 277
x"01350",-- 309
x"01350",-- 309
x"010e0",-- 270
x"00b10",-- 177
x"00140",-- 20
x"ff6d0",-- -147
x"fec80",-- -312
x"fe5f0",-- -417
x"fe390",-- -455
x"fe280",-- -472
x"fe2d0",-- -467
x"fe160",-- -490
x"fe080",-- -504
x"fdf30",-- -525
x"fdf60",-- -522
x"fe490",-- -439
x"feb70",-- -329
x"ff310",-- -207
x"ffc10",-- -63
x"005c0",-- 92
x"00dc0",-- 220
x"013b0",-- 315
x"01880",-- 392
x"01990",-- 409
x"01b30",-- 435
x"01b30",-- 435
x"01940",-- 404
x"01650",-- 357
x"01120",-- 274
x"00870",-- 135
x"ffea0",-- -22
x"ff860",-- -122
x"ff510",-- -175
x"ff0c0",-- -244
x"fead0",-- -339
x"fe7f0",-- -385
x"fea20",-- -350
x"feb90",-- -327
x"fecd0",-- -307
x"fede0",-- -290
x"ff070",-- -249
x"ff2b0",-- -213
x"ff4e0",-- -178
x"ff8b0",-- -117
x"ffc40",-- -60
x"00080",-- 8
x"00260",-- 38
x"00670",-- 103
x"00a70",-- 167
x"00bb0",-- 187
x"00c10",-- 193
x"00aa0",-- 170
x"00b10",-- 177
x"00b60",-- 182
x"00de0",-- 222
x"00e10",-- 225
x"00c60",-- 198
x"00c80",-- 200
x"00cf0",-- 207
x"00d20",-- 210
x"00cf0",-- 207
x"00930",-- 147
x"00410",-- 65
x"fff80",-- -8
x"ffbc0",-- -68
x"ff920",-- -110
x"ff790",-- -135
x"ff5d0",-- -163
x"ff380",-- -200
x"ff3f0",-- -193
x"ff4e0",-- -178
x"ff650",-- -155
x"ff630",-- -157
x"ff5e0",-- -162
x"ff7c0",-- -132
x"ffdf0",-- -33
x"00500",-- 80
x"00b90",-- 185
x"010b0",-- 267
x"01450",-- 325
x"01800",-- 384
x"018a0",-- 394
x"01600",-- 352
x"01290",-- 297
x"00e10",-- 225
x"00940",-- 148
x"005d0",-- 93
x"00300",-- 48
x"fff90",-- -7
x"ff990",-- -103
x"ff380",-- -200
x"fedf0",-- -289
x"fea20",-- -350
x"fea50",-- -347
x"febe0",-- -322
x"fed50",-- -299
x"ff020",-- -254
x"ff420",-- -190
x"ff9c0",-- -100
x"ffe70",-- -25
x"00170",-- 23
x"00410",-- 65
x"005d0",-- 93
x"00760",-- 118
x"00a00",-- 160
x"00e10",-- 225
x"00fa0",-- 250
x"01090",-- 265
x"00dc0",-- 220
x"00800",-- 128
x"002f0",-- 47
x"ffc40",-- -60
x"ff800",-- -128
x"ff4c0",-- -180
x"ff300",-- -208
x"ff440",-- -188
x"ff4f0",-- -177
x"ff600",-- -160
x"ff510",-- -175
x"ff4f0",-- -177
x"ff6c0",-- -148
x"ff970",-- -105
x"ffdd0",-- -35
x"000f0",-- 15
x"00490",-- 73
x"00870",-- 135
x"00990",-- 153
x"00890",-- 137
x"00570",-- 87
x"00280",-- 40
x"00030",-- 3
x"00020",-- 2
x"001b0",-- 27
x"002b0",-- 43
x"00430",-- 67
x"00570",-- 87
x"00700",-- 112
x"006b0",-- 107
x"006e0",-- 110
x"00570",-- 87
x"00530",-- 83
x"00570",-- 87
x"003c0",-- 60
x"00260",-- 38
x"00070",-- 7
x"ffdf0",-- -33
x"ffb00",-- -80
x"ff880",-- -120
x"ff740",-- -140
x"ff630",-- -157
x"ff5d0",-- -163
x"ff630",-- -157
x"ff680",-- -152
x"ff710",-- -143
x"ff830",-- -125
x"ff990",-- -103
x"ffb80",-- -72
x"ffef0",-- -17
x"00160",-- 22
x"003f0",-- 63
x"005a0",-- 90
x"00620",-- 98
x"006b0",-- 107
x"006c0",-- 108
x"00500",-- 80
x"003c0",-- 60
x"002b0",-- 43
x"00200",-- 32
x"00120",-- 18
x"ffee0",-- -18
x"ffad0",-- -83
x"ff670",-- -153
x"ff310",-- -207
x"ff0e0",-- -242
x"ff040",-- -252
x"ff070",-- -249
x"ff070",-- -249
x"ff220",-- -222
x"ff510",-- -175
x"ff790",-- -135
x"ffb70",-- -73
x"fff40",-- -12
x"00110",-- 17
x"000a0",-- 10
x"00020",-- 2
x"00050",-- 5
x"001b0",-- 27
x"00160",-- 22
x"00120",-- 18
x"00140",-- 20
x"00110",-- 17
x"00210",-- 33
x"000c0",-- 12
x"00050",-- 5
x"ffec0",-- -20
x"ffdd0",-- -35
x"ffe00",-- -32
x"ffef0",-- -17
x"ffea0",-- -22
x"ffd10",-- -47
x"ffc90",-- -55
x"ffb50",-- -75
x"ffb80",-- -72
x"ffa40",-- -92
x"ffa30",-- -93
x"ffa60",-- -90
x"ffab0",-- -85
x"ffbc0",-- -68
x"ffbc0",-- -68
x"ffbf0",-- -65
x"ffb80",-- -72
x"ffc60",-- -58
x"ffda0",-- -38
x"fffb0",-- -5
x"001b0",-- 27
x"003c0",-- 60
x"005f0",-- 95
x"00820",-- 130
x"009e0",-- 158
x"009d0",-- 157
x"008e0",-- 142
x"006c0",-- 108
x"004e0",-- 78
x"00370",-- 55
x"001c0",-- 28
x"fffe0",-- -2
x"fff80",-- -8
x"ffe20",-- -30
x"ffc90",-- -55
x"ffa60",-- -90
x"ff970",-- -105
x"ffa30",-- -93
x"ff9c0",-- -100
x"ffb50",-- -75
x"ffdd0",-- -35
x"00050",-- 5
x"00280",-- 40
x"003e0",-- 62
x"00530",-- 83
x"005d0",-- 93
x"00640",-- 100
x"007a0",-- 122
x"008e0",-- 142
x"00870",-- 135
x"00840",-- 132
x"00730",-- 115
x"005a0",-- 90
x"003a0",-- 58
x"00030",-- 3
x"ffd50",-- -43
x"ffbf0",-- -65
x"ffb00",-- -80
x"ffba0",-- -70
x"ffda0",-- -38
x"ffdb0",-- -37
x"ffe90",-- -23
x"ffec0",-- -20
x"00020",-- 2
x"000f0",-- 15
x"00280",-- 40
x"004e0",-- 78
x"00760",-- 118
x"00ad0",-- 173
x"00b70",-- 183
x"00bc0",-- 188
x"00960",-- 150
x"00610",-- 97
x"00350",-- 53
x"00280",-- 40
x"00170",-- 23
x"00160",-- 22
x"001c0",-- 28
x"00110",-- 17
x"001b0",-- 27
x"00160",-- 22
x"00050",-- 5
x"00050",-- 5
x"00000",-- 0
x"00170",-- 23
x"00300",-- 48
x"002a0",-- 42
x"00160",-- 22
x"000a0",-- 10
x"fffe0",-- -2
x"ffe00",-- -32
x"ffe50",-- -27
x"ffea0",-- -22
x"fff40",-- -12
x"fffe0",-- -2
x"00000",-- 0
x"fffe0",-- -2
x"00000",-- 0
x"fffb0",-- -5
x"fff10",-- -15
x"00000",-- 0
x"000c0",-- 12
x"00210",-- 33
x"00350",-- 53
x"00530",-- 83
x"00440",-- 68
x"002d0",-- 45
x"00160",-- 22
x"fff90",-- -7
x"ffdd0",-- -35
x"ffcb0",-- -53
x"ffda0",-- -38
x"ffda0",-- -38
x"ffd10",-- -47
x"ffd50",-- -43
x"ffc20",-- -62
x"ffae0",-- -82
x"ffa80",-- -88
x"ff9c0",-- -100
x"ff9a0",-- -102
x"ffa10",-- -95
x"ffdb0",-- -37
x"fffe0",-- -2
x"00120",-- 18
x"002f0",-- 47
x"002f0",-- 47
x"00410",-- 65
x"00460",-- 70
x"00480",-- 72
x"00340",-- 52
x"000c0",-- 12
x"fff80",-- -8
x"ffe40",-- -28
x"ffea0",-- -22
x"ffea0",-- -22
x"ffdb0",-- -37
x"ffc70",-- -57
x"ffba0",-- -70
x"ffc40",-- -60
x"ffc20",-- -62
x"ffb80",-- -72
x"ffa90",-- -87
x"ffb70",-- -73
x"ffd50",-- -43
x"ffe50",-- -27
x"ffea0",-- -22
x"ffdd0",-- -35
x"ffd10",-- -47
x"ffd00",-- -48
x"ffd80",-- -40
x"ffe50",-- -27
x"ffd50",-- -43
x"ffdb0",-- -37
x"ffda0",-- -38
x"ffea0",-- -22
x"fff90",-- -7
x"fff40",-- -12
x"fff90",-- -7
x"fff80",-- -8
x"00020",-- 2
x"00000",-- 0
x"00050",-- 5
x"00080",-- 8
x"00050",-- 5
x"000c0",-- 12
x"00080",-- 8
x"00080",-- 8
x"00000",-- 0
x"ffdf0",-- -33
x"ffce0",-- -50
x"ffbd0",-- -67
x"ffba0",-- -70
x"ffb20",-- -78
x"ffb70",-- -73
x"ffc20",-- -62
x"ffbf0",-- -65
x"ffd50",-- -43
x"fff10",-- -15
x"00000",-- 0
x"000c0",-- 12
x"000f0",-- 15
x"00170",-- 23
x"00230",-- 35
x"002b0",-- 43
x"002b0",-- 43
x"002b0",-- 43
x"00280",-- 40
x"001c0",-- 28
x"000f0",-- 15
x"00020",-- 2
x"fffe0",-- -2
x"fff60",-- -10
x"ffdb0",-- -37
x"ffc60",-- -58
x"ffbc0",-- -68
x"ffb80",-- -72
x"ffc90",-- -55
x"ffc10",-- -63
x"ffc60",-- -58
x"ffd30",-- -45
x"ffe70",-- -25
x"fffe0",-- -2
x"000f0",-- 15
x"00250",-- 37
x"003c0",-- 60
x"00570",-- 87
x"004e0",-- 78
x"00460",-- 70
x"003a0",-- 58
x"00370",-- 55
x"003a0",-- 58
x"001e0",-- 30
x"00020",-- 2
x"ffea0",-- -22
x"ffcc0",-- -52
x"ffbf0",-- -65
x"ffb80",-- -72
x"ffbc0",-- -68
x"ffb50",-- -75
x"ffc90",-- -55
x"ffda0",-- -38
x"fff10",-- -15
x"00050",-- 5
x"000f0",-- 15
x"001b0",-- 27
x"00210",-- 33
x"00200",-- 32
x"00110",-- 17
x"00110",-- 17
x"00000",-- 0
x"00080",-- 8
x"fffe0",-- -2
x"ffe70",-- -25
x"ffe40",-- -28
x"ffdb0",-- -37
x"ffdd0",-- -35
x"ffd10",-- -47
x"ffd10",-- -47
x"ffd50",-- -43
x"ffe20",-- -30
x"ffe50",-- -27
x"ffee0",-- -18
x"fffb0",-- -5
x"00030",-- 3
x"000c0",-- 12
x"fffe0",-- -2
x"00000",-- 0
x"00020",-- 2
x"fff80",-- -8
x"fff60",-- -10
x"fff80",-- -8
x"fffd0",-- -3
x"fff10",-- -15
x"fff40",-- -12
x"fff80",-- -8
x"fff30",-- -13
x"fff10",-- -15
x"fff60",-- -10
x"fffe0",-- -2
x"00000",-- 0
x"fffb0",-- -5
x"fffb0",-- -5
x"00030",-- 3
x"00160",-- 22
x"00210",-- 33
x"00200",-- 32
x"002f0",-- 47
x"00210",-- 33
x"001e0",-- 30
x"00160",-- 22
x"00080",-- 8
x"fffe0",-- -2
x"ffdf0",-- -33
x"ffd10",-- -47
x"ffd30",-- -45
x"ffe70",-- -25
x"fff10",-- -15
x"fff10",-- -15
x"ffea0",-- -22
x"ffec0",-- -20
x"ffee0",-- -18
x"ffe00",-- -32
x"ffe70",-- -25
x"ffea0",-- -22
x"fffb0",-- -5
x"00250",-- 37
x"00350",-- 53
x"002a0",-- 42
x"001b0",-- 27
x"000f0",-- 15
x"000f0",-- 15
x"00000",-- 0
x"fffb0",-- -5
x"fff80",-- -8
x"000a0",-- 10
x"00280",-- 40
x"002b0",-- 43
x"00250",-- 37
x"000a0",-- 10
x"fffe0",-- -2
x"000a0",-- 10
x"00030",-- 3
x"00000",-- 0
x"00140",-- 20
x"00020",-- 2
x"ffd80",-- -40
x"ffd00",-- -48
x"ffee0",-- -18
x"ffef0",-- -17
x"fffd0",-- -3
x"00020",-- 2
x"00000",-- 0
x"000f0",-- 15
x"00280",-- 40
x"00170",-- 23
x"ffda0",-- -38
x"ffe90",-- -23
x"fff80",-- -8
x"00160",-- 22
x"003e0",-- 62
x"00480",-- 72
x"00620",-- 98
x"00690",-- 105
x"00760",-- 118
x"00760",-- 118
x"005a0",-- 90
x"00460",-- 70
x"003c0",-- 60
x"002f0",-- 47
x"002f0",-- 47
x"00320",-- 50
x"00390",-- 57
x"002a0",-- 42
x"00170",-- 23
x"00080",-- 8
x"000a0",-- 10
x"00200",-- 32
x"001c0",-- 28
x"00260",-- 38
x"003f0",-- 63
x"004b0",-- 75
x"004b0",-- 75
x"003c0",-- 60
x"00340",-- 52
x"001e0",-- 30
x"001b0",-- 27
x"00210",-- 33
x"00200",-- 32
x"001b0",-- 27
x"001c0",-- 28
x"00030",-- 3
x"fff80",-- -8
x"fff40",-- -12
x"ffdf0",-- -33
x"ffd10",-- -47
x"ffd10",-- -47
x"ffdf0",-- -33
x"fff60",-- -10
x"00000",-- 0
x"000c0",-- 12
x"00080",-- 8
x"00050",-- 5
x"00080",-- 8
x"00120",-- 18
x"00160",-- 22
x"00160",-- 22
x"001e0",-- 30
x"00110",-- 17
x"000f0",-- 15
x"00080",-- 8
x"fffd0",-- -3
x"fff40",-- -12
x"fff80",-- -8
x"ffe90",-- -23
x"fff40",-- -12
x"fffd0",-- -3
x"00050",-- 5
x"00080",-- 8
x"fff10",-- -15
x"fff60",-- -10
x"ffee0",-- -18
x"ffe50",-- -27
x"fff30",-- -13
x"00020",-- 2
x"000a0",-- 10
x"fffd0",-- -3
x"fffb0",-- -5
x"fff10",-- -15
x"ffe50",-- -27
x"ffdb0",-- -37
x"ffd30",-- -45
x"ffad0",-- -83
x"ff970",-- -105
x"ffc10",-- -63
x"ffdf0",-- -33
x"ffe50",-- -27
x"ffd80",-- -40
x"ffce0",-- -50
x"ffc90",-- -55
x"ffc60",-- -58
x"ffce0",-- -50
x"ffdb0",-- -37
x"ffd60",-- -42
x"ffdb0",-- -37
x"ffe70",-- -25
x"fff40",-- -12
x"fff40",-- -12
x"ffe50",-- -27
x"ffe20",-- -30
x"ffdf0",-- -33
x"ffdd0",-- -35
x"ffe50",-- -27
x"ffe00",-- -32
x"ffcc0",-- -52
x"ffbc0",-- -68
x"ffb50",-- -75
x"ffc20",-- -62
x"ffd80",-- -40
x"ffb50",-- -75
x"ff8a0",-- -118
x"ff830",-- -125
x"ffb00",-- -80
x"ffc20",-- -62
x"ffba0",-- -70
x"ffb20",-- -78
x"ffbc0",-- -68
x"ffbd0",-- -67
x"ffa90",-- -87
x"ffc90",-- -55
x"ffb70",-- -73
x"ffb80",-- -72
x"ffbf0",-- -65
x"ffcb0",-- -53
x"ffce0",-- -50
x"ffbd0",-- -67
x"ffb80",-- -72
x"ff670",-- -153
x"ff3b0",-- -197
x"ff9e0",-- -98
x"ffda0",-- -38
x"fff40",-- -12
x"00070",-- 7
x"fff80",-- -8
x"ffdf0",-- -33
x"ffe20",-- -30
x"ffc90",-- -55
x"ffae0",-- -82
x"ffc20",-- -62
x"ffc40",-- -60
x"ffe40",-- -28
x"00110",-- 17
x"00190",-- 25
x"000d0",-- 13
x"00120",-- 18
x"001b0",-- 27
x"000f0",-- 15
x"001b0",-- 27
x"00300",-- 48
x"002b0",-- 43
x"00300",-- 48
x"00320",-- 50
x"003a0",-- 58
x"003a0",-- 58
x"001c0",-- 28
x"00000",-- 0
x"00000",-- 0
x"001c0",-- 28
x"00210",-- 33
x"00000",-- 0
x"ffe50",-- -27
x"ffd30",-- -45
x"ffea0",-- -22
x"ffea0",-- -22
x"fff40",-- -12
x"00000",-- 0
x"fff90",-- -7
x"ffef0",-- -17
x"ffe20",-- -30
x"000f0",-- 15
x"00080",-- 8
x"000a0",-- 10
x"00000",-- 0
x"ffee0",-- -18
x"ffdd0",-- -35
x"ffea0",-- -22
x"fff90",-- -7
x"ffe90",-- -23
x"ffec0",-- -20
x"ffe20",-- -30
x"ffe40",-- -28
x"fff10",-- -15
x"ffea0",-- -22
x"ffe40",-- -28
x"ffea0",-- -22
x"ffdf0",-- -33
x"ffe50",-- -27
x"fff10",-- -15
x"00050",-- 5
x"fff40",-- -12
x"fff40",-- -12
x"00000",-- 0
x"00030",-- 3
x"fffb0",-- -5
x"00000",-- 0
x"00190",-- 25
x"000c0",-- 12
x"00140",-- 20
x"00050",-- 5
x"fffb0",-- -5
x"fff40",-- -12
x"ffe50",-- -27
x"ffd60",-- -42
x"ffe40",-- -28
x"00000",-- 0
x"ffee0",-- -18
x"fff40",-- -12
x"fff80",-- -8
x"fff10",-- -15
x"00000",-- 0
x"ffee0",-- -18
x"00080",-- 8
x"00080",-- 8
x"00050",-- 5
x"000a0",-- 10
x"000f0",-- 15
x"000f0",-- 15
x"fffe0",-- -2
x"fff40",-- -12
x"fff60",-- -10
x"fff80",-- -8
x"ffdb0",-- -37
x"fff10",-- -15
x"fffb0",-- -5
x"ffe20",-- -30
x"fff40",-- -12
x"00020",-- 2
x"fff90",-- -7
x"fffe0",-- -2
x"000c0",-- 12
x"00020",-- 2
x"fff40",-- -12
x"00020",-- 2
x"00120",-- 18
x"fff90",-- -7
x"fffe0",-- -2
x"ffe90",-- -23
x"fff60",-- -10
x"000a0",-- 10
x"fffb0",-- -5
x"fff40",-- -12
x"ffe50",-- -27
x"ffd50",-- -43
x"ffd10",-- -47
x"ffd00",-- -48
x"fff80",-- -8
x"00160",-- 22
x"fffb0",-- -5
x"00110",-- 17
x"00250",-- 37
x"001b0",-- 27
x"000f0",-- 15
x"ffef0",-- -17
x"ffe50",-- -27
x"ffd00",-- -48
x"fff80",-- -8
x"fffe0",-- -2
x"fffb0",-- -5
x"00080",-- 8
x"fff90",-- -7
x"fffb0",-- -5
x"fff30",-- -13
x"ffd50",-- -43
x"ffc60",-- -58
x"ffb30",-- -77
x"ffd30",-- -45
x"ffe00",-- -32
x"ffd50",-- -43
x"ffdb0",-- -37
x"ffd80",-- -40
x"ffcb0",-- -53
x"ffb80",-- -72
x"ffd50",-- -43
x"fff40",-- -12
x"fff60",-- -10
x"ffe20",-- -30
x"ffd10",-- -47
x"ffd00",-- -48
x"ffe40",-- -28
x"ffd30",-- -45
x"ff9e0",-- -98
x"ff950",-- -107
x"ff9f0",-- -97
x"ffb20",-- -78
x"ffb30",-- -77
x"ff990",-- -103
x"ffa90",-- -87
x"ff8f0",-- -113
x"ff600",-- -160
x"ff9a0",-- -102
x"ffa30",-- -93
x"ff970",-- -105
x"ffc60",-- -58
x"ffad0",-- -83
x"ffcb0",-- -53
x"ffd30",-- -45
x"ffa30",-- -93
x"ffa60",-- -90
x"ff8d0",-- -115
x"ffa90",-- -87
x"ff9f0",-- -97
x"ffa90",-- -87
x"ffdd0",-- -35
x"ffb80",-- -72
x"ffbc0",-- -68
x"ffcb0",-- -53
x"ffd30",-- -45
x"ffc90",-- -55
x"ff990",-- -103
x"ff830",-- -125
x"ff8a0",-- -118
x"ffc10",-- -63
x"ffee0",-- -18
x"ffb00",-- -80
x"ffa40",-- -92
x"ffa90",-- -87
x"ff800",-- -128
x"ffbc0",-- -68
x"ff9f0",-- -97
x"ff990",-- -103
x"ffd10",-- -47
x"ff900",-- -112
x"ffd10",-- -47
x"fffb0",-- -5
x"ffab0",-- -85
x"ffa10",-- -95
x"ffa90",-- -87
x"ff9c0",-- -100
x"ffc70",-- -57
x"ffd10",-- -47
x"ffc60",-- -58
x"ffe40",-- -28
x"ffef0",-- -17
x"ffba0",-- -70
x"000c0",-- 12
x"ffe40",-- -28
x"ffa60",-- -90
x"ffdf0",-- -33
x"fff10",-- -15
x"00000",-- 0
x"ffa30",-- -93
x"ffce0",-- -50
x"ffab0",-- -85
x"ff9f0",-- -97
x"ffb80",-- -72
x"ff810",-- -127
x"ff7b0",-- -133
x"ff810",-- -127
x"ff580",-- -168
x"ff970",-- -105
x"00080",-- 8
x"fffe0",-- -2
x"000f0",-- 15
x"ffee0",-- -18
x"ffe50",-- -27
x"00170",-- 23
x"00000",-- 0
x"ffec0",-- -20
x"ffea0",-- -22
x"004b0",-- 75
x"00280",-- 40
x"00050",-- 5
x"00490",-- 73
x"00280",-- 40
x"00320",-- 50
x"00430",-- 67
x"00660",-- 102
x"00520",-- 82
x"ffd50",-- -43
x"005a0",-- 90
x"008a0",-- 138
x"00030",-- 3
x"00530",-- 83
x"fff10",-- -15
x"ffb50",-- -75
x"00000",-- 0
x"ffd10",-- -47
x"ffa30",-- -93
x"ffe20",-- -30
x"00030",-- 3
x"ffe00",-- -32
x"00190",-- 25
x"005a0",-- 90
x"00430",-- 67
x"ffda0",-- -38
x"fffb0",-- -5
x"000d0",-- 13
x"00080",-- 8
x"fff40",-- -12
x"000a0",-- 10
x"005d0",-- 93
x"fffb0",-- -5
x"00750",-- 117
x"000c0",-- 12
x"00080",-- 8
x"00a80",-- 168
x"00320",-- 50
x"003a0",-- 58
x"00960",-- 150
x"00990",-- 153
x"fff30",-- -13
x"00370",-- 55
x"00610",-- 97
x"ffef0",-- -17
x"00120",-- 18
x"00580",-- 88
x"00990",-- 153
x"003c0",-- 60
x"ffcb0",-- -53
x"00690",-- 105
x"00320",-- 50
x"ffc60",-- -58
x"00440",-- 68
x"00a80",-- 168
x"00520",-- 82
x"00200",-- 32
x"00f00",-- 240
x"01150",-- 277
x"003c0",-- 60
x"000d0",-- 13
x"00a00",-- 160
x"ffdd0",-- -35
x"ffd50",-- -43
x"00b10",-- 177
x"ffe70",-- -25
x"00570",-- 87
x"014f0",-- 335
x"00b60",-- 182
x"00700",-- 112
x"00840",-- 132
x"004d0",-- 77
x"ffc40",-- -60
x"00870",-- 135
x"003a0",-- 58
x"ffbc0",-- -68
x"003e0",-- 62
x"00b20",-- 178
x"ffc40",-- -60
x"00850",-- 133
x"01880",-- 392
x"00430",-- 67
x"00a80",-- 168
x"003e0",-- 62
x"ff4a0",-- -182
x"fed20",-- -302
x"fee40",-- -284
x"00430",-- 67
x"01e50",-- 485
x"006e0",-- 110
x"ffd80",-- -40
x"01490",-- 329
x"010e0",-- 270
x"01470",-- 327
x"fe120",-- -494
x"fdf30",-- -525
x"ff990",-- -103
x"02ad0",-- 685
x"01380",-- 312
x"01bf0",-- 447
x"036c0",-- 876
x"fd130",-- -749
x"ff4e0",-- -178
x"01270",-- 295
x"fec10",-- -319
x"fd470",-- -697
x"009d0",-- 157
x"026b0",-- 619
x"005d0",-- 93
x"02c60",-- 710
x"00020",-- 2
x"fd290",-- -727
x"ff970",-- -105
x"ffe40",-- -28
x"ff2e0",-- -210
x"ff060",-- -250
x"00a00",-- 160
x"ffb00",-- -80
x"00670",-- 103
x"03210",-- 801
x"02210",-- 545
x"fd680",-- -664
x"fd790",-- -647
x"025f0",-- 607
x"02ff0",-- 767
x"fff60",-- -10
x"00a50",-- 165
x"016d0",-- 365
x"fd680",-- -664
x"ffc20",-- -62
x"02980",-- 664
x"ff380",-- -200
x"fdda0",-- -550
x"00f40",-- 244
x"feb20",-- -334
x"ff100",-- -240
x"04300",-- 1072
x"ffb50",-- -75
x"fe2d0",-- -467
x"021c0",-- 540
x"011a0",-- 282
x"00eb0",-- 235
x"00230",-- 35
x"ff5b0",-- -165
x"fe3a0",-- -454
x"fde90",-- -535
x"fdbc0",-- -580
x"ffdb0",-- -37
x"00da0",-- 218
x"fc8f0",-- -881
x"01770",-- 375
x"00640",-- 100
x"fcc30",-- -829
x"00a80",-- 168
x"fc070",-- -1017
x"fc6c0",-- -916
x"febb0",-- -325
x"ff450",-- -187
x"01e50",-- 485
x"00d40",-- 212
x"ffc20",-- -62
x"fc7a0",-- -902
x"02d90",-- 729
x"03120",-- 786
x"fe9d0",-- -355
x"01b20",-- 434
x"003c0",-- 60
x"ff470",-- -185
x"042a0",-- 1066
x"03760",-- 886
x"02480",-- 584
x"01ec0",-- 492
x"00d90",-- 217
x"02530",-- 595
x"00050",-- 5
x"01c60",-- 454
x"ffb20",-- -78
x"ffee0",-- -18
x"00620",-- 98
x"00480",-- 72
x"01cc0",-- 460
x"fdf10",-- -527
x"fe1e0",-- -482
x"fea80",-- -344
x"fddf0",-- -545
x"01710",-- 369
x"ff900",-- -112
x"fde40",-- -540
x"01bd0",-- 445
x"01470",-- 327
x"01d60",-- 470
x"01dd0",-- 477
x"ff6a0",-- -150
x"00ad0",-- 173
x"00f90",-- 249
x"00a80",-- 168
x"02ea0",-- 746
x"02f00",-- 752
x"01260",-- 294
x"ff260",-- -218
x"04f50",-- 1269
x"04820",-- 1154
x"fe700",-- -400
x"01ad0",-- 429
x"02af0",-- 687
x"00e80",-- 232
x"01a60",-- 422
x"02c60",-- 710
x"00eb0",-- 235
x"fe8a0",-- -374
x"fe960",-- -362
x"01f60",-- 502
x"00080",-- 8
x"fe620",-- -414
x"005a0",-- 90
x"fe300",-- -464
x"01c70",-- 455
x"044b0",-- 1099
x"00000",-- 0
x"fec10",-- -319
x"ff6a0",-- -150
x"00df0",-- 223
x"ffee0",-- -18
x"00160",-- 22
x"019e0",-- 414
x"ffa40",-- -92
x"ff800",-- -128
x"006b0",-- 107
x"00460",-- 70
x"ff850",-- -123
x"fe410",-- -447
x"00f90",-- 249
x"ff1d0",-- -227
x"fe3a0",-- -454
x"019e0",-- 414
x"02120",-- 530
x"ff5b0",-- -165
x"fea20",-- -350
x"02cd0",-- 717
x"02c30",-- 707
x"031c0",-- 796
x"ffef0",-- -17
x"fc2b0",-- -981
x"00930",-- 147
x"008a0",-- 138
x"ff620",-- -158
x"02300",-- 560
x"fd3b0",-- -709
x"fe890",-- -375
x"01220",-- 290
x"fe390",-- -455
x"ffee0",-- -18
x"01040",-- 260
x"009d0",-- 157
x"fe070",-- -505
x"000c0",-- 12
x"fe050",-- -507
x"ff4a0",-- -182
x"01830",-- 387
x"fc840",-- -892
x"fefa0",-- -262
x"00df0",-- 223
x"ff680",-- -152
x"00050",-- 5
x"ffe90",-- -23
x"00500",-- 80
x"fec50",-- -315
x"fe1e0",-- -482
x"02210",-- 545
x"fd3f0",-- -705
x"001b0",-- 27
x"00d50",-- 213
x"ff830",-- -125
x"ff7c0",-- -132
x"fe7b0",-- -389
x"fea70",-- -345
x"fc9e0",-- -866
x"fefc0",-- -260
x"fd7c0",-- -644
x"fda40",-- -604
x"003a0",-- 58
x"026e0",-- 622
x"feaa0",-- -342
x"fed70",-- -297
x"03300",-- 816
x"fe070",-- -505
x"fe140",-- -492
x"fe050",-- -507
x"fe2f0",-- -465
x"ff590",-- -167
x"ff290",-- -215
x"00570",-- 87
x"fe210",-- -479
x"01350",-- 309
x"fe700",-- -400
x"ff240",-- -220
x"00dc0",-- 220
x"fc1c0",-- -996
x"fe7a0",-- -390
x"00490",-- 73
x"fd9c0",-- -612
x"01580",-- 344
x"fe6e0",-- -402
x"fe350",-- -459
x"020a0",-- 522
x"fdd00",-- -560
x"ff560",-- -170
x"ffc90",-- -55
x"ffbf0",-- -65
x"ffc20",-- -62
x"002d0",-- 45
x"ffd10",-- -47
x"ff5e0",-- -162
x"01300",-- 304
x"ff310",-- -207
x"ff4a0",-- -182
x"ffd00",-- -48
x"ffc70",-- -57
x"01810",-- 385
x"ffee0",-- -18
x"ff110",-- -239
x"fdfb0",-- -517
x"ff150",-- -235
x"fdae0",-- -594
x"fe930",-- -365
x"00200",-- 32
x"feeb0",-- -277
x"ffea0",-- -22
x"ff440",-- -188
x"fe7b0",-- -389
x"015e0",-- 350
x"fe530",-- -429
x"ff830",-- -125
x"ff6a0",-- -150
x"fd530",-- -685
x"007d0",-- 125
x"fda80",-- -600
x"fff80",-- -8
x"01d30",-- 467
x"fe070",-- -505
x"00020",-- 2
x"fda10",-- -607
x"fe6e0",-- -402
x"ffea0",-- -22
x"fdbc0",-- -580
x"01f30",-- 499
x"fe800",-- -384
x"ff9e0",-- -98
x"ff590",-- -167
x"01130",-- 275
x"00730",-- 115
x"fe190",-- -487
x"01a90",-- 425
x"fd060",-- -762
x"00a70",-- 167
x"ffc20",-- -62
x"fe8e0",-- -370
x"03ea0",-- 1002
x"fdec0",-- -532
x"011f0",-- 287
x"01b30",-- 435
x"fde70",-- -537
x"02030",-- 515
x"fde00",-- -544
x"ff4c0",-- -180
x"014c0",-- 332
x"ff6a0",-- -150
x"fdea0",-- -534
x"ff360",-- -202
x"00c80",-- 200
x"fe620",-- -414
x"01e20",-- 482
x"00a00",-- 160
x"00df0",-- 223
x"ff740",-- -140
x"fe6b0",-- -405
x"002f0",-- 47
x"00700",-- 112
x"00440",-- 68
x"02460",-- 582
x"00e10",-- 225
x"00640",-- 100
x"02460",-- 582
x"ff630",-- -157
x"02750",-- 629
x"ff150",-- -235
x"00a20",-- 162
x"01b00",-- 432
x"ffb00",-- -80
x"00640",-- 100
x"00e80",-- 232
x"feed0",-- -275
x"00b10",-- 177
x"fc550",-- -939
x"022f0",-- 559
x"00ef0",-- 239
x"fd720",-- -654
x"04ea0",-- 1258
x"fbd60",-- -1066
x"036c0",-- 876
x"fdda0",-- -550
x"00a20",-- 162
x"ffce0",-- -50
x"00140",-- 20
x"00d90",-- 217
x"01220",-- 290
x"01e20",-- 482
x"fc300",-- -976
x"01d10",-- 465
x"009b0",-- 155
x"fff40",-- -12
x"ffbf0",-- -65
x"ff940",-- -108
x"ff060",-- -250
x"03860",-- 902
x"fe000",-- -512
x"00610",-- 97
x"ffc60",-- -58
x"fcb70",-- -841
x"01f60",-- 502
x"fe4d0",-- -435
x"fdda0",-- -550
x"020c0",-- 524
x"fed70",-- -297
x"00e40",-- 228
x"018d0",-- 397
x"fd240",-- -732
x"ff8f0",-- -113
x"008e0",-- 142
x"fc520",-- -942
x"00520",-- 82
x"02e00",-- 736
x"01360",-- 310
x"01670",-- 359
x"fde00",-- -544
x"020d0",-- 525
x"ff450",-- -187
x"00230",-- 35
x"008e0",-- 142
x"fe570",-- -425
x"02930",-- 659
x"ff1a0",-- -230
x"fe8f0",-- -369
x"00960",-- 150
x"ffee0",-- -18
x"fed90",-- -295
x"00a20",-- 162
x"004e0",-- 78
x"fe460",-- -442
x"ff800",-- -128
x"ffdf0",-- -33
x"ff7e0",-- -130
x"00840",-- 132
x"fd670",-- -665
x"00f50",-- 245
x"ff9e0",-- -98
x"fe610",-- -415
x"01290",-- 297
x"feb40",-- -332
x"00d20",-- 210
x"fdda0",-- -550
x"023f0",-- 575
x"fee60",-- -282
x"00730",-- 115
x"ffda0",-- -38
x"fe5f0",-- -417
x"02e00",-- 736
x"fab70",-- -1353
x"00bb0",-- 187
x"ff4a0",-- -182
x"fc940",-- -876
x"027f0",-- 639
x"fd1b0",-- -741
x"ffc70",-- -57
x"015b0",-- 347
x"fdc10",-- -575
x"01cc0",-- 460
x"ffe20",-- -30
x"ff260",-- -218
x"ff3a0",-- -198
x"000f0",-- 15
x"00020",-- 2
x"ff9f0",-- -97
x"00440",-- 68
x"ff9c0",-- -100
x"00f50",-- 245
x"ff970",-- -105
x"01030",-- 259
x"00d90",-- 217
x"fe620",-- -414
x"002a0",-- 42
x"00c50",-- 197
x"fe9b0",-- -357
x"01100",-- 272
x"ff130",-- -237
x"fe340",-- -460
x"00f20",-- 242
x"fec10",-- -319
x"ffd00",-- -48
x"ff9e0",-- -98
x"fe440",-- -444
x"01450",-- 325
x"ff090",-- -247
x"ff540",-- -172
x"004e0",-- 78
x"fe820",-- -382
x"01650",-- 357
x"000c0",-- 12
x"00710",-- 113
x"00cb0",-- 203
x"00440",-- 68
x"fe3a0",-- -454
x"00ed0",-- 237
x"ffa30",-- -93
x"ff990",-- -103
x"01ad0",-- 429
x"fe250",-- -475
x"008f0",-- 143
x"ff070",-- -249
x"ffc10",-- -63
x"016f0",-- 367
x"024b0",-- 587
x"ffd80",-- -40
x"00b90",-- 185
x"ff800",-- -128
x"fd920",-- -622
x"00af0",-- 175
x"ff350",-- -203
x"ffc10",-- -63
x"ff210",-- -223
x"00340",-- 52
x"ff8d0",-- -115
x"01d50",-- 469
x"ffd10",-- -47
x"000d0",-- 13
x"002b0",-- 43
x"ff8a0",-- -118
x"00a80",-- 168
x"fe520",-- -430
x"ffe50",-- -27
x"fe6c0",-- -404
x"00c30",-- 195
x"00710",-- 113
x"00cb0",-- 203
x"ff830",-- -125
x"ff510",-- -175
x"01010",-- 257
x"fec50",-- -315
x"00640",-- 100
x"001b0",-- 27
x"00280",-- 40
x"00f00",-- 240
x"feff0",-- -257
x"ffbd0",-- -67
x"fee80",-- -280
x"014e0",-- 334
x"ff800",-- -128
x"00e80",-- 232
x"ffbc0",-- -68
x"00b60",-- 182
x"023e0",-- 574
x"00000",-- 0
x"01f90",-- 505
x"ff5b0",-- -165
x"011f0",-- 287
x"fea80",-- -344
x"00d50",-- 213
x"ff800",-- -128
x"fefa0",-- -262
x"00160",-- 22
x"ff3b0",-- -197
x"01c20",-- 450
x"001b0",-- 27
x"00cf0",-- 207
x"ff5d0",-- -163
x"ffc10",-- -63
x"ff790",-- -135
x"ff600",-- -160
x"ff5e0",-- -162
x"00260",-- 38
x"00080",-- 8
x"00020",-- 2
x"ffe70",-- -25
x"ff3a0",-- -198
x"01710",-- 369
x"00410",-- 65
x"031d0",-- 797
x"01810",-- 385
x"00a70",-- 167
x"01600",-- 352
x"febc0",-- -324
x"01170",-- 279
x"ff0e0",-- -242
x"ff740",-- -140
x"008c0",-- 140
x"00e80",-- 232
x"00d00",-- 208
x"015d0",-- 349
x"ff0e0",-- -242
x"ff6a0",-- -150
x"001b0",-- 27
x"ff440",-- -188
x"01d30",-- 467
x"ffdb0",-- -37
x"00670",-- 103
x"015e0",-- 350
x"fed20",-- -302
x"00b90",-- 185
x"003a0",-- 58
x"003a0",-- 58
x"ff8b0",-- -117
x"00000",-- 0
x"00b60",-- 182
x"001e0",-- 30
x"022d0",-- 557
x"ff6a0",-- -150
x"01400",-- 320
x"001b0",-- 27
x"ff790",-- -135
x"ffbf0",-- -65
x"ff900",-- -112
x"fdf10",-- -527
x"ffb00",-- -80
x"ff350",-- -203
x"fe890",-- -375
x"00550",-- 85
x"00640",-- 100
x"01030",-- 259
x"01e20",-- 482
x"002d0",-- 45
x"00a30",-- 163
x"00f90",-- 249
x"fff80",-- -8
x"00120",-- 18
x"ffec0",-- -20
x"ff760",-- -138
x"00210",-- 33
x"ffec0",-- -20
x"009d0",-- 157
x"01ae0",-- 430
x"00940",-- 148
x"00ff0",-- 255
x"ff6d0",-- -147
x"ff800",-- -128
x"ff3f0",-- -193
x"00a80",-- 168
x"ffc20",-- -62
x"01310",-- 305
x"fe9b0",-- -357
x"feb20",-- -334
x"007b0",-- 123
x"fe820",-- -382
x"ffe70",-- -25
x"fe6e0",-- -402
x"ffa30",-- -93
x"ff850",-- -123
x"008e0",-- 142
x"00620",-- 98
x"ff720",-- -142
x"019e0",-- 414
x"ffb80",-- -72
x"00660",-- 102
x"fef00",-- -272
x"fdf80",-- -520
x"00a70",-- 167
x"fe7b0",-- -389
x"00390",-- 57
x"00c60",-- 198
x"ff0c0",-- -244
x"00f50",-- 245
x"ffdf0",-- -33
x"ffb20",-- -78
x"005d0",-- 93
x"ff620",-- -158
x"006e0",-- 110
x"00050",-- 5
x"002f0",-- 47
x"ff540",-- -172
x"ff350",-- -203
x"ffc90",-- -55
x"00350",-- 53
x"008c0",-- 140
x"011a0",-- 282
x"fff40",-- -12
x"fff30",-- -13
x"00440",-- 68
x"ffc90",-- -55
x"00300",-- 48
x"ff4f0",-- -177
x"00d70",-- 215
x"ff940",-- -108
x"ffb80",-- -72
x"ffb20",-- -78
x"feda0",-- -294
x"ff110",-- -239
x"fe730",-- -397
x"ff670",-- -153
x"ff6f0",-- -145
x"ffc70",-- -57
x"00c50",-- 197
x"ff8f0",-- -113
x"00120",-- 18
x"01300",-- 304
x"ff4e0",-- -178
x"002b0",-- 43
x"ffb30",-- -77
x"fee60",-- -282
x"ff860",-- -122
x"ff710",-- -143
x"00030",-- 3
x"008f0",-- 143
x"00b60",-- 182
x"000f0",-- 15
x"008c0",-- 140
x"ff4a0",-- -182
x"00bc0",-- 188
x"00640",-- 100
x"00670",-- 103
x"00f90",-- 249
x"00390",-- 57
x"feb10",-- -335
x"ff5b0",-- -165
x"ff4e0",-- -178
x"ffa60",-- -90
x"00430",-- 67
x"fe9e0",-- -354
x"003a0",-- 58
x"ff4a0",-- -182
x"ff8b0",-- -117
x"01080",-- 264
x"ff810",-- -127
x"ffe40",-- -28
x"fef00",-- -272
x"001c0",-- 28
x"feb90",-- -327
x"fef00",-- -272
x"00690",-- 105
x"fe670",-- -409
x"01b30",-- 435
x"ff210",-- -223
x"01740",-- 372
x"ff5e0",-- -162
x"00280",-- 40
x"00a00",-- 160
x"ff490",-- -183
x"028a0",-- 650
x"fe0d0",-- -499
x"01560",-- 342
x"fed50",-- -299
x"00370",-- 55
x"00dc0",-- 220
x"ff7c0",-- -132
x"00480",-- 72
x"fff40",-- -12
x"006e0",-- 110
x"00480",-- 72
x"005c0",-- 92
x"ff630",-- -157
x"ff800",-- -128
x"ff620",-- -158
x"ffe00",-- -32
x"ff990",-- -103
x"fec80",-- -312
x"fed70",-- -297
x"ff540",-- -172
x"005c0",-- 92
x"ff1a0",-- -230
x"000c0",-- 12
x"00000",-- 0
x"ff0b0",-- -245
x"00b10",-- 177
x"ffb20",-- -78
x"00cf0",-- 207
x"ff510",-- -175
x"ffe00",-- -32
x"ffe20",-- -30
x"ffb80",-- -72
x"ffec0",-- -20
x"ffce0",-- -50
x"00160",-- 22
x"ffdb0",-- -37
x"fffb0",-- -5
x"00350",-- 53
x"00ca0",-- 202
x"ffc20",-- -62
x"00ef0",-- 239
x"ffdb0",-- -37
x"fff30",-- -13
x"ffef0",-- -17
x"ffa10",-- -95
x"ffbf0",-- -65
x"ff100",-- -240
x"003a0",-- 58
x"ffa90",-- -87
x"00050",-- 5
x"00800",-- 128
x"fe800",-- -384
x"ffea0",-- -22
x"ffad0",-- -83
x"ffa60",-- -90
x"00d90",-- 217
x"00120",-- 18
x"003e0",-- 62
x"ff2e0",-- -210
x"00570",-- 87
x"febc0",-- -324
x"00280",-- 40
x"ffe50",-- -27
x"fe320",-- -462
x"00620",-- 98
x"fee40",-- -284
x"ff630",-- -157
x"001b0",-- 27
x"ff110",-- -239
x"00a80",-- 168
x"ffe50",-- -27
x"ffda0",-- -38
x"ffc20",-- -62
x"00140",-- 20
x"001e0",-- 30
x"003f0",-- 63
x"ff3b0",-- -197
x"fff40",-- -12
x"ffad0",-- -83
x"00a80",-- 168
x"001b0",-- 27
x"fff40",-- -12
x"fff90",-- -7
x"ffb80",-- -72
x"008f0",-- 143
x"ffe40",-- -28
x"00b10",-- 177
x"ffad0",-- -83
x"001e0",-- 30
x"fe190",-- -487
x"00050",-- 5
x"ffb30",-- -77
x"ffe20",-- -30
x"005d0",-- 93
x"00070",-- 7
x"00410",-- 65
x"ffce0",-- -50
x"003a0",-- 58
x"fe690",-- -407
x"00b90",-- 185
x"ff710",-- -143
x"ff580",-- -168
x"00020",-- 2
x"ff580",-- -168
x"004d0",-- 77
x"003c0",-- 60
x"ffdb0",-- -37
x"ffa60",-- -90
x"00ac0",-- 172
x"fef70",-- -265
x"00210",-- 33
x"00000",-- 0
x"002b0",-- 43
x"01c90",-- 457
x"00850",-- 133
x"00f00",-- 240
x"010b0",-- 267
x"ff210",-- -223
x"ff2e0",-- -210
x"003a0",-- 58
x"fe5d0",-- -419
x"004e0",-- 78
x"ff070",-- -249
x"ffb30",-- -77
x"000f0",-- 15
x"00440",-- 68
x"ff860",-- -122
x"ffc90",-- -55
x"ff8f0",-- -113
x"fe5d0",-- -419
x"00000",-- 0
x"ff310",-- -207
x"00210",-- 33
x"008e0",-- 142
x"00c50",-- 197
x"00190",-- 25
x"00d20",-- 210
x"ff6a0",-- -150
x"ffef0",-- -17
x"01220",-- 290
x"ff670",-- -153
x"00ac0",-- 172
x"ff240",-- -220
x"00670",-- 103
x"010d0",-- 269
x"fe610",-- -415
x"008c0",-- 140
x"feac0",-- -340
x"00a30",-- 163
x"ff800",-- -128
x"fe990",-- -359
x"00aa0",-- 170
x"feaf0",-- -337
x"014e0",-- 334
x"ff310",-- -207
x"00410",-- 65
x"ff950",-- -107
x"00120",-- 18
x"01210",-- 289
x"ff040",-- -252
x"015b0",-- 347
x"fff90",-- -7
x"00730",-- 115
x"013f0",-- 319
x"00620",-- 98
x"003e0",-- 62
x"016d0",-- 365
x"fef20",-- -270
x"ff950",-- -107
x"00340",-- 52
x"ffee0",-- -18
x"00070",-- 7
x"ffba0",-- -70
x"ff380",-- -200
x"ffc90",-- -55
x"00050",-- 5
x"feb90",-- -327
x"ff0b0",-- -245
x"ff3b0",-- -197
x"ffd60",-- -42
x"ff740",-- -140
x"ffe00",-- -32
x"fffe0",-- -2
x"00000",-- 0
x"00800",-- 128
x"01040",-- 260
x"00250",-- 37
x"ff9e0",-- -98
x"ffe00",-- -32
x"ff150",-- -235
x"007d0",-- 125
x"ffc10",-- -63
x"01ef0",-- 495
x"02480",-- 584
x"00000",-- 0
x"03970",-- 919
x"ff6d0",-- -147
x"01560",-- 342
x"00ad0",-- 173
x"fea20",-- -350
x"014e0",-- 334
x"feb90",-- -327
x"00500",-- 80
x"ffd30",-- -45
x"ff240",-- -220
x"fff80",-- -8
x"ff270",-- -217
x"01100",-- 272
x"fe2a0",-- -470
x"ff310",-- -207
x"ff710",-- -143
x"fdbc0",-- -580
x"000d0",-- 13
x"fe7d0",-- -387
x"fff10",-- -15
x"ff2e0",-- -210
x"00500",-- 80
x"ffce0",-- -50
x"00120",-- 18
x"019a0",-- 410
x"fef30",-- -269
x"01dd0",-- 477
x"00d70",-- 215
x"00800",-- 128
x"007d0",-- 125
x"fecd0",-- -307
x"006b0",-- 107
x"ff7c0",-- -132
x"ffc60",-- -58
x"01060",-- 262
x"ff9c0",-- -100
x"003e0",-- 62
x"00df0",-- 223
x"00a80",-- 168
x"00170",-- 23
x"ffc40",-- -60
x"ffda0",-- -38
x"ffdf0",-- -33
x"005c0",-- 92
x"000c0",-- 12
x"00980",-- 152
x"002f0",-- 47
x"ffae0",-- -82
x"ff900",-- -112
x"00f20",-- 242
x"00490",-- 73
x"00050",-- 5
x"004d0",-- 77
x"fea80",-- -344
x"00710",-- 113
x"00750",-- 117
x"00550",-- 85
x"ffb20",-- -78
x"ffe00",-- -32
x"01970",-- 407
x"fec30",-- -317
x"ffe20",-- -30
x"ff6a0",-- -150
x"00390",-- 57
x"00960",-- 150
x"00000",-- 0
x"01010",-- 257
x"ff8b0",-- -117
x"00430",-- 67
x"ff760",-- -138
x"003c0",-- 60
x"00700",-- 112
x"ff110",-- -239
x"00700",-- 112
x"006e0",-- 110
x"ffe20",-- -30
x"016a0",-- 362
x"fef50",-- -267
x"ff860",-- -122
x"00c00",-- 192
x"ff5b0",-- -165
x"01900",-- 400
x"003a0",-- 58
x"ffd80",-- -40
x"011c0",-- 284
x"ffda0",-- -38
x"00660",-- 102
x"00a30",-- 163
x"feac0",-- -340
x"014f0",-- 335
x"ffe00",-- -32
x"00820",-- 130
x"022b0",-- 555
x"ff380",-- -200
x"00e10",-- 225
x"ff830",-- -125
x"00050",-- 5
x"ffd50",-- -43
x"ff7c0",-- -132
x"ff790",-- -135
x"ff1f0",-- -225
x"010d0",-- 269
x"fe910",-- -367
x"ff2b0",-- -213
x"ff630",-- -157
x"ff1c0",-- -228
x"01290",-- 297
x"fec30",-- -317
x"ffec0",-- -20
x"00390",-- 57
x"ff6a0",-- -150
x"003c0",-- 60
x"ffb80",-- -72
x"ff990",-- -103
x"013b0",-- 315
x"ffa60",-- -90
x"01c60",-- 454
x"003f0",-- 63
x"007a0",-- 122
x"00f00",-- 240
x"ffbc0",-- -68
x"01030",-- 259
x"ff6c0",-- -148
x"02930",-- 659
x"ff110",-- -239
x"01790",-- 377
x"ffdf0",-- -33
x"ff600",-- -160
x"01450",-- 325
x"fd8b0",-- -629
x"002f0",-- 47
x"fe930",-- -365
x"ff6d0",-- -147
x"00190",-- 25
x"ff900",-- -112
x"00530",-- 83
x"ff800",-- -128
x"00b20",-- 178
x"fef70",-- -265
x"015e0",-- 350
x"ffd00",-- -48
x"ffce0",-- -50
x"01770",-- 375
x"febb0",-- -325
x"01380",-- 312
x"00350",-- 53
x"ff940",-- -108
x"005d0",-- 93
x"009b0",-- 155
x"01060",-- 262
x"012b0",-- 299
x"002f0",-- 47
x"ffd80",-- -40
x"fff10",-- -15
x"ff9c0",-- -100
x"ff760",-- -138
x"ff4f0",-- -177
x"ff7b0",-- -133
x"ff6a0",-- -150
x"00480",-- 72
x"ff210",-- -223
x"00370",-- 55
x"00b20",-- 178
x"ff510",-- -175
x"012c0",-- 300
x"fffe0",-- -2
x"00640",-- 100
x"01900",-- 400
x"ff6a0",-- -150
x"002a0",-- 42
x"ffc20",-- -62
x"ffbd0",-- -67
x"00dc0",-- 220
x"ff560",-- -170
x"008c0",-- 140
x"013b0",-- 315
x"fff80",-- -8
x"01c10",-- 449
x"ff470",-- -185
x"ffdf0",-- -33
x"ff7c0",-- -132
x"ffa30",-- -93
x"00000",-- 0
x"006b0",-- 107
x"003f0",-- 63
x"fe850",-- -379
x"014e0",-- 334
x"fed20",-- -302
x"ff800",-- -128
x"fef00",-- -272
x"fee60",-- -282
x"ffea0",-- -22
x"00dc0",-- 220
x"fff10",-- -15
x"ffec0",-- -20
x"ffd00",-- -48
x"00800",-- 128
x"00c00",-- 192
x"ffbc0",-- -68
x"ff760",-- -138
x"010d0",-- 269
x"00280",-- 40
x"015e0",-- 350
x"01310",-- 305
x"fe460",-- -442
x"00fe0",-- 254
x"ff180",-- -232
x"01e00",-- 480
x"003e0",-- 62
x"00000",-- 0
x"00020",-- 2
x"ffd60",-- -42
x"ffd50",-- -43
x"00550",-- 85
x"ffb00",-- -80
x"ff5d0",-- -163
x"ff900",-- -112
x"00840",-- 132
x"005c0",-- 92
x"feee0",-- -274
x"ffe50",-- -27
x"fe570",-- -425
x"00c50",-- 197
x"fe8f0",-- -369
x"ffee0",-- -18
x"00120",-- 18
x"ff470",-- -185
x"01560",-- 342
x"00110",-- 17
x"00b90",-- 185
x"002b0",-- 43
x"fee40",-- -284
x"00b90",-- 185
x"002b0",-- 43
x"ffc20",-- -62
x"01580",-- 344
x"fede0",-- -290
x"01060",-- 262
x"00bb0",-- 187
x"00340",-- 52
x"01350",-- 309
x"ff6a0",-- -150
x"fff10",-- -15
x"ffe50",-- -27
x"fffb0",-- -5
x"00230",-- 35
x"ffda0",-- -38
x"ffce0",-- -50
x"ff880",-- -120
x"00da0",-- 218
x"fff10",-- -15
x"fe620",-- -414
x"00d20",-- 210
x"feaf0",-- -337
x"015b0",-- 347
x"ffbf0",-- -65
x"ffbd0",-- -67
x"01380",-- 312
x"fe6b0",-- -405
x"01da0",-- 474
x"fdf80",-- -520
x"018a0",-- 394
x"ff130",-- -237
x"ff9f0",-- -97
x"01900",-- 400
x"ff2c0",-- -212
x"01df0",-- 479
x"ff240",-- -220
x"00930",-- 147
x"ffc40",-- -60
x"003e0",-- 62
x"00700",-- 112
x"ff670",-- -153
x"ffa90",-- -87
x"ff830",-- -125
x"febb0",-- -325
x"011f0",-- 287
x"ffdb0",-- -37
x"ff850",-- -123
x"00a50",-- 165
x"fe710",-- -399
x"00840",-- 132
x"ffee0",-- -18
x"00f50",-- 245
x"fef30",-- -269
x"016c0",-- 364
x"fffe0",-- -2
x"ff580",-- -168
x"006b0",-- 107
x"fe3e0",-- -450
x"00f20",-- 242
x"00050",-- 5
x"00530",-- 83
x"00120",-- 18
x"ffec0",-- -20
x"ff5e0",-- -162
x"ff510",-- -175
x"00440",-- 68
x"ff040",-- -252
x"003a0",-- 58
x"ff770",-- -137
x"00af0",-- 175
x"002b0",-- 43
x"00fe0",-- 254
x"ffa90",-- -87
x"00710",-- 113
x"ff8d0",-- -115
x"ff540",-- -172
x"01060",-- 262
x"ffad0",-- -83
x"ff710",-- -143
x"ffe20",-- -30
x"00530",-- 83
x"ff180",-- -232
x"01360",-- 310
x"fead0",-- -339
x"006b0",-- 107
x"fede0",-- -290
x"ff7c0",-- -132
x"ff270",-- -217
x"fea80",-- -344
x"00410",-- 65
x"ff950",-- -107
x"00b20",-- 178
x"001e0",-- 30
x"ff770",-- -137
x"00690",-- 105
x"ff7c0",-- -132
x"01a60",-- 422
x"ffe40",-- -28
x"00410",-- 65
x"ffc70",-- -57
x"ff210",-- -223
x"fffb0",-- -5
x"ffd50",-- -43
x"011a0",-- 282
x"fe6c0",-- -404
x"01360",-- 310
x"009e0",-- 158
x"015e0",-- 350
x"00850",-- 133
x"002a0",-- 42
x"fedf0",-- -289
x"ff6d0",-- -147
x"ff5d0",-- -163
x"ff070",-- -249
x"011f0",-- 287
x"fedf0",-- -289
x"00410",-- 65
x"fead0",-- -339
x"fffd0",-- -3
x"ff600",-- -160
x"fee40",-- -284
x"013d0",-- 317
x"ff4f0",-- -177
x"01490",-- 329
x"fec50",-- -315
x"feda0",-- -294
x"ffdf0",-- -33
x"000c0",-- 12
x"01380",-- 312
x"ffe90",-- -23
x"ffe90",-- -23
x"00b60",-- 182
x"00730",-- 115
x"ffdb0",-- -37
x"00250",-- 37
x"ff6c0",-- -148
x"00730",-- 115
x"00120",-- 18
x"00c10",-- 193
x"00460",-- 70
x"00440",-- 68
x"ffe50",-- -27
x"ff810",-- -127
x"01150",-- 277
x"fed40",-- -300
x"ff1c0",-- -228
x"fe3e0",-- -450
x"ffc20",-- -62
x"00940",-- 148
x"ff8d0",-- -115
x"00b10",-- 177
x"00340",-- 52
x"ff090",-- -247
x"003c0",-- 60
x"fda30",-- -605
x"ff920",-- -110
x"ff6a0",-- -150
x"ff7c0",-- -132
x"01950",-- 405
x"fffe0",-- -2
x"032e0",-- 814
x"ffcc0",-- -52
x"00690",-- 105
x"fedf0",-- -289
x"008c0",-- 140
x"ff950",-- -107
x"ff4c0",-- -180
x"007b0",-- 123
x"fef30",-- -269
x"00370",-- 55
x"ff850",-- -123
x"ff6a0",-- -150
x"ff110",-- -239
x"ff420",-- -190
x"fff90",-- -7
x"fe3e0",-- -450
x"ff1c0",-- -228
x"ff470",-- -185
x"fe280",-- -472
x"ffa90",-- -87
x"ff530",-- -173
x"01170",-- 279
x"00080",-- 8
x"00480",-- 72
x"ffc60",-- -58
x"02b70",-- 695
x"018a0",-- 394
x"00390",-- 57
x"ffdd0",-- -35
x"fe9d0",-- -355
x"00980",-- 152
x"ff950",-- -107
x"feed0",-- -275
x"00a30",-- 163
x"00160",-- 22
x"002b0",-- 43
x"02000",-- 512
x"ff380",-- -200
x"01210",-- 289
x"ff770",-- -137
x"fea80",-- -344
x"ffa30",-- -93
x"fde40",-- -540
x"ff0e0",-- -242
x"ffa80",-- -88
x"00570",-- 87
x"00210",-- 33
x"00b40",-- 180
x"008c0",-- 140
x"ffd30",-- -45
x"00b60",-- 182
x"002a0",-- 42
x"ff0c0",-- -244
x"fff60",-- -10
x"fe9d0",-- -355
x"fef30",-- -269
x"00610",-- 97
x"feeb0",-- -277
x"00b20",-- 178
x"ff950",-- -107
x"ff4a0",-- -182
x"00200",-- 32
x"ff4f0",-- -177
x"ffab0",-- -85
x"fec30",-- -317
x"01670",-- 359
x"ffd10",-- -47
x"ffe50",-- -27
x"00d20",-- 210
x"00b90",-- 185
x"016d0",-- 365
x"ffa90",-- -87
x"fff30",-- -13
x"ff540",-- -172
x"ff740",-- -140
x"ffa10",-- -95
x"00c00",-- 192
x"00280",-- 40
x"fecd0",-- -307
x"00dc0",-- 220
x"ff9f0",-- -97
x"fe370",-- -457
x"ff0c0",-- -244
x"fe1b0",-- -485
x"00f70",-- 247
x"00670",-- 103
x"00530",-- 83
x"02ad0",-- 685
x"ffb80",-- -72
x"01150",-- 277
x"ff010",-- -255
x"00ad0",-- 173
x"fe730",-- -397
x"ffd80",-- -40
x"02f40",-- 756
x"fe200",-- -480
x"02980",-- 664
x"009d0",-- 157
x"00c50",-- 197
x"ffa30",-- -93
x"fd7c0",-- -644
x"fff10",-- -15
x"fe940",-- -364
x"01ad0",-- 429
x"feff0",-- -257
x"fef20",-- -270
x"00dc0",-- 220
x"fef00",-- -272
x"00320",-- 50
x"fe340",-- -460
x"ff150",-- -235
x"01240",-- 292
x"ff830",-- -125
x"00020",-- 2
x"013a0",-- 314
x"00d20",-- 210
x"005f0",-- 95
x"ffdb0",-- -37
x"fefa0",-- -262
x"ff040",-- -252
x"02ad0",-- 685
x"00580",-- 88
x"01310",-- 305
x"01fe0",-- 510
x"ffc10",-- -63
x"02030",-- 515
x"ff1c0",-- -228
x"00140",-- 20
x"011c0",-- 284
x"fe870",-- -377
x"00990",-- 153
x"002f0",-- 47
x"fedf0",-- -289
x"00640",-- 100
x"feaf0",-- -337
x"ff740",-- -140
x"ff3a0",-- -198
x"ffa60",-- -90
x"fea70",-- -345
x"ff6a0",-- -150
x"00c60",-- 198
x"fe0f0",-- -497
x"01a60",-- 422
x"feeb0",-- -277
x"fe750",-- -395
x"014e0",-- 334
x"01030",-- 259
x"00ff0",-- 255
x"fefc0",-- -260
x"003c0",-- 60
x"00a30",-- 163
x"ff790",-- -135
x"00a50",-- 165
x"00c50",-- 197
x"00b90",-- 185
x"ff850",-- -123
x"00b20",-- 178
x"00480",-- 72
x"01920",-- 402
x"00260",-- 38
x"fe020",-- -510
x"00ef0",-- 239
x"00b20",-- 178
x"fe460",-- -442
x"00020",-- 2
x"ff630",-- -157
x"fed90",-- -295
x"016a0",-- 362
x"ff800",-- -128
x"00b10",-- 177
x"ff580",-- -168
x"01120",-- 274
x"01e20",-- 482
x"01650",-- 357
x"ff5e0",-- -162
x"fe530",-- -429
x"00960",-- 150
x"fefc0",-- -260
x"00490",-- 73
x"fe550",-- -427
x"ffc90",-- -55
x"01130",-- 275
x"002f0",-- 47
x"013b0",-- 315
x"ffd50",-- -43
x"ff5d0",-- -163
x"ff380",-- -200
x"00730",-- 115
x"fef50",-- -267
x"fe0f0",-- -497
x"fe9e0",-- -354
x"00850",-- 133
x"00840",-- 132
x"ff470",-- -185
x"036c0",-- 876
x"00e80",-- 232
x"01490",-- 329
x"ff800",-- -128
x"00b70",-- 183
x"00120",-- 18
x"ff510",-- -175
x"00610",-- 97
x"00af0",-- 175
x"029e0",-- 670
x"ff740",-- -140
x"00e30",-- 227
x"00080",-- 8
x"fec50",-- -315
x"00260",-- 38
x"fe8a0",-- -374
x"ff6a0",-- -150
x"ffdb0",-- -37
x"018a0",-- 394
x"01c10",-- 449
x"fede0",-- -290
x"fec60",-- -314
x"feeb0",-- -277
x"ff6a0",-- -150
x"ff3a0",-- -198
x"fef20",-- -270
x"ff680",-- -152
x"ff790",-- -135
x"00c30",-- 195
x"001b0",-- 27
x"00cb0",-- 203
x"00c50",-- 197
x"00080",-- 8
x"02070",-- 519
x"00230",-- 35
x"01ef0",-- 495
x"00120",-- 18
x"ffce0",-- -50
x"014c0",-- 332
x"ffea0",-- -22
x"01fe0",-- 510
x"005a0",-- 90
x"008f0",-- 143
x"00d90",-- 217
x"01360",-- 310
x"02370",-- 567
x"fecf0",-- -305
x"ff9c0",-- -100
x"ff240",-- -220
x"ff2e0",-- -210
x"001c0",-- 28
x"fe7d0",-- -387
x"00ef0",-- 239
x"ff100",-- -240
x"ff420",-- -190
x"00660",-- 102
x"ff800",-- -128
x"fde50",-- -539
x"fdb00",-- -592
x"00c80",-- 200
x"00000",-- 0
x"00e60",-- 230
x"02020",-- 514
x"00e90",-- 233
x"01cc0",-- 460
x"01260",-- 294
x"00af0",-- 175
x"01b80",-- 440
x"003f0",-- 63
x"01950",-- 405
x"00ac0",-- 172
x"ffbd0",-- -67
x"fede0",-- -290
x"00980",-- 152
x"ffc70",-- -57
x"fd630",-- -669
x"fdc10",-- -575
x"fe930",-- -365
x"00250",-- 37
x"ff270",-- -217
x"00440",-- 68
x"015e0",-- 350
x"01650",-- 357
x"ffd50",-- -43
x"ff670",-- -153
x"ff540",-- -172
x"ff450",-- -187
x"fffe0",-- -2
x"003e0",-- 62
x"007a0",-- 122
x"01860",-- 390
x"01c70",-- 455
x"005f0",-- 95
x"02020",-- 514
x"ffdd0",-- -35
x"00610",-- 97
x"008f0",-- 143
x"fe9b0",-- -357
x"00500",-- 80
x"00250",-- 37
x"00870",-- 135
x"fffe0",-- -2
x"001b0",-- 27
x"febb0",-- -325
x"002a0",-- 42
x"00800",-- 128
x"003e0",-- 62
x"009e0",-- 158
x"ff880",-- -120
x"ff3b0",-- -197
x"fe870",-- -377
x"00750",-- 117
x"ffa30",-- -93
x"00000",-- 0
x"00910",-- 145
x"016d0",-- 365
x"017c0",-- 380
x"01630",-- 355
x"00430",-- 67
x"ffc70",-- -57
x"ff420",-- -190
x"fef00",-- -272
x"00710",-- 113
x"ffb20",-- -78
x"ff020",-- -254
x"ff8d0",-- -115
x"01c90",-- 457
x"01120",-- 274
x"00530",-- 83
x"ff3b0",-- -197
x"00840",-- 132
x"ffd60",-- -42
x"00d00",-- 208
x"01e20",-- 482
x"ff540",-- -172
x"00480",-- 72
x"004e0",-- 78
x"00430",-- 67
x"01650",-- 357
x"fe570",-- -425
x"00ef0",-- 239
x"01260",-- 294
x"ff3f0",-- -193
x"ff920",-- -110
x"ff6a0",-- -150
x"01060",-- 262
x"00530",-- 83
x"ffa40",-- -92
x"ff670",-- -153
x"ffa90",-- -87
x"fe8e0",-- -370
x"fe6e0",-- -402
x"011f0",-- 287
x"015e0",-- 350
x"ff9f0",-- -97
x"02350",-- 565
x"00320",-- 50
x"01180",-- 280
x"ffdb0",-- -37
x"fee10",-- -287
x"ff3a0",-- -198
x"fdef0",-- -529
x"01860",-- 390
x"000f0",-- 15
x"fd5d0",-- -675
x"ff380",-- -200
x"ffb20",-- -78
x"01ec0",-- 492
x"ff650",-- -155
x"fefa0",-- -262
x"01f10",-- 497
x"016c0",-- 364
x"02000",-- 512
x"ff7e0",-- -130
x"fea20",-- -350
x"fdd10",-- -559
x"ffc40",-- -60
x"00440",-- 68
x"ff580",-- -168
x"01260",-- 294
x"ff950",-- -107
x"00930",-- 147
x"03ae0",-- 942
x"fe890",-- -375
x"003e0",-- 62
x"ffb50",-- -75
x"fe250",-- -475
x"00fc0",-- 252
x"fe210",-- -479
x"fee10",-- -287
x"fe550",-- -427
x"fe9d0",-- -355
x"ffd60",-- -42
x"00000",-- 0
x"002f0",-- 47
x"fef00",-- -272
x"01040",-- 260
x"01d80",-- 472
x"00930",-- 147
x"00070",-- 7
x"fef00",-- -272
x"ff1d0",-- -227
x"ff540",-- -172
x"fe530",-- -429
x"01290",-- 297
x"ff450",-- -187
x"01580",-- 344
x"014e0",-- 334
x"00670",-- 103
x"01540",-- 340
x"fe800",-- -384
x"00c00",-- 192
x"ff5e0",-- -162
x"fecd0",-- -307
x"fe350",-- -459
x"ff790",-- -135
x"ff5e0",-- -162
x"fefc0",-- -260
x"ffa60",-- -90
x"fde70",-- -537
x"ffc20",-- -62
x"ff9c0",-- -100
x"fff90",-- -7
x"00f90",-- 249
x"ff7b0",-- -133
x"ffba0",-- -70
x"00b10",-- 177
x"ffa80",-- -88
x"ffb50",-- -75
x"00d40",-- 212
x"00760",-- 118
x"015b0",-- 347
x"00d70",-- 215
x"ffa30",-- -93
x"01090",-- 265
x"ffbc0",-- -68
x"fd9e0",-- -610
x"fd770",-- -649
x"ff600",-- -160
x"ff310",-- -207
x"ffd60",-- -42
x"ff360",-- -202
x"00160",-- 22
x"01830",-- 387
x"ff580",-- -168
x"ff220",-- -222
x"fe280",-- -472
x"ffc60",-- -58
x"013a0",-- 314
x"00820",-- 130
x"00000",-- 0
x"ffa30",-- -93
x"00120",-- 18
x"01b00",-- 432
x"00070",-- 7
x"ff400",-- -192
x"005a0",-- 90
x"ffbd0",-- -67
x"00280",-- 40
x"011a0",-- 282
x"ffef0",-- -17
x"fff40",-- -12
x"006e0",-- 110
x"fd4e0",-- -690
x"ff9c0",-- -100
x"ff620",-- -158
x"ff1a0",-- -230
x"ff990",-- -103
x"fcfd0",-- -771
x"00640",-- 100
x"01e70",-- 487
x"021e0",-- 542
x"ffce0",-- -50
x"ffa30",-- -93
x"ffbc0",-- -68
x"00b90",-- 185
x"00320",-- 50
x"008c0",-- 140
x"00210",-- 33
x"00c00",-- 192
x"008f0",-- 143
x"00140",-- 20
x"00e60",-- 230
x"fd560",-- -682
x"00bc0",-- 188
x"fddf0",-- -545
x"ff8d0",-- -115
x"03210",-- 801
x"fdd50",-- -555
x"ffd30",-- -45
x"ffad0",-- -83
x"00120",-- 18
x"01d10",-- 465
x"fe6c0",-- -404
x"fe640",-- -412
x"fffb0",-- -5
x"ff9c0",-- -100
x"ff940",-- -108
x"01b70",-- 439
x"001e0",-- 30
x"fe7f0",-- -385
x"02930",-- 659
x"00620",-- 98
x"00e40",-- 228
x"02460",-- 582
x"fdcc0",-- -564
x"02110",-- 529
x"004d0",-- 77
x"ff880",-- -120
x"027f0",-- 639
x"fdb30",-- -589
x"fdfe0",-- -514
x"ff8d0",-- -115
x"fee40",-- -284
x"00930",-- 147
x"ff380",-- -200
x"fed40",-- -300
x"00dc0",-- 220
x"ff9f0",-- -97
x"ffe70",-- -25
x"00730",-- 115
x"00500",-- 80
x"00a80",-- 168
x"00480",-- 72
x"01330",-- 307
x"00aa0",-- 170
x"007f0",-- 127
x"ff210",-- -223
x"ffdb0",-- -37
x"fe820",-- -382
x"ff6d0",-- -147
x"00930",-- 147
x"00ff0",-- 255
x"01260",-- 294
x"01310",-- 305
x"00cf0",-- 207
x"00410",-- 65
x"ffba0",-- -70
x"fe3a0",-- -454
x"ffce0",-- -50
x"ff6c0",-- -148
x"00440",-- 68
x"00f20",-- 242
x"feb10",-- -335
x"fe690",-- -407
x"ff0b0",-- -245
x"ffd10",-- -47
x"004e0",-- 78
x"ff790",-- -135
x"ffd50",-- -43
x"001e0",-- 30
x"ffa10",-- -95
x"00c60",-- 198
x"ffe00",-- -32
x"fef00",-- -272
x"ff8a0",-- -118
x"002b0",-- 43
x"ffb20",-- -78
x"00730",-- 115
x"00530",-- 83
x"00020",-- 2
x"00980",-- 152
x"00000",-- 0
x"006e0",-- 110
x"ffce0",-- -50
x"001b0",-- 27
x"00210",-- 33
x"00c00",-- 192
x"02d70",-- 727
x"fea30",-- -349
x"01130",-- 275
x"ff650",-- -155
x"fe350",-- -459
x"00660",-- 102
x"fe140",-- -492
x"00840",-- 132
x"fed70",-- -297
x"ff6d0",-- -147
x"013b0",-- 315
x"ff860",-- -122
x"ff990",-- -103
x"00430",-- 67
x"fe7d0",-- -387
x"ff0e0",-- -242
x"00730",-- 115
x"00610",-- 97
x"00d20",-- 210
x"008c0",-- 140
x"ffa90",-- -87
x"01ba0",-- 442
x"ff580",-- -168
x"00050",-- 5
x"ffec0",-- -20
x"fe3a0",-- -454
x"fff40",-- -12
x"018b0",-- 395
x"004b0",-- 75
x"01380",-- 312
x"ff800",-- -128
x"006c0",-- 108
x"01030",-- 259
x"00f50",-- 245
x"ff5d0",-- -163
x"fe3e0",-- -450
x"01170",-- 279
x"ff740",-- -140
x"00d00",-- 208
x"00840",-- 132
x"fe2d0",-- -467
x"ff2b0",-- -213
x"fde00",-- -544
x"ff4e0",-- -178
x"00c60",-- 198
x"fe480",-- -440
x"00c00",-- 192
x"ff8a0",-- -118
x"00530",-- 83
x"fea80",-- -344
x"00dc0",-- 220
x"ff010",-- -255
x"fe6b0",-- -405
x"02160",-- 534
x"00a30",-- 163
x"01270",-- 295
x"ff970",-- -105
x"01c10",-- 449
x"011a0",-- 282
x"ffd80",-- -40
x"00230",-- 35
x"00550",-- 85
x"fff10",-- -15
x"00000",-- 0
x"00f20",-- 242
x"00550",-- 85
x"00a80",-- 168
x"ff6d0",-- -147
x"00820",-- 130
x"ff270",-- -217
x"fe7a0",-- -390
x"ff440",-- -188
x"ff9c0",-- -100
x"ff5d0",-- -163
x"ffc40",-- -60
x"ffdb0",-- -37
x"003e0",-- 62
x"01b70",-- 439
x"ff800",-- -128
x"ffcb0",-- -53
x"004d0",-- 77
x"ffb20",-- -78
x"01130",-- 275
x"00df0",-- 223
x"00c50",-- 197
x"003c0",-- 60
x"ff800",-- -128
x"00280",-- 40
x"ff9c0",-- -100
x"00730",-- 115
x"00700",-- 112
x"01d30",-- 467
x"00160",-- 22
x"fff40",-- -12
x"01170",-- 279
x"00c10",-- 193
x"ffa30",-- -93
x"ff0e0",-- -242
x"ff800",-- -128
x"ff9c0",-- -100
x"011f0",-- 287
x"00210",-- 33
x"fec50",-- -315
x"000a0",-- 10
x"01b70",-- 439
x"007a0",-- 122
x"00fc0",-- 252
x"ff100",-- -240
x"00000",-- 0
x"005a0",-- 90
x"00050",-- 5
x"00660",-- 102
x"ffc90",-- -55
x"00580",-- 88
x"00370",-- 55
x"ffba0",-- -70
x"ff9c0",-- -100
x"ff400",-- -192
x"ff0e0",-- -242
x"007a0",-- 122
x"00160",-- 22
x"00480",-- 72
x"00d50",-- 213
x"00c80",-- 200
x"00a00",-- 160
x"00990",-- 153
x"00410",-- 65
x"feff0",-- -257
x"fea80",-- -344
x"000c0",-- 12
x"ffbd0",-- -67
x"00280",-- 40
x"01180",-- 280
x"01030",-- 259
x"00a00",-- 160
x"00300",-- 48
x"00bc0",-- 188
x"ffbf0",-- -65
x"009d0",-- 157
x"008e0",-- 142
x"ff540",-- -172
x"00be0",-- 190
x"ffda0",-- -38
x"ffa30",-- -93
x"00670",-- 103
x"00670",-- 103
x"ffa10",-- -95
x"ff420",-- -190
x"ff630",-- -157
x"00480",-- 72
x"003c0",-- 60
x"ffb70",-- -73
x"ff1d0",-- -227
x"00440",-- 68
x"00800",-- 128
x"ff070",-- -249
x"013b0",-- 315
x"ff3f0",-- -193
x"00250",-- 37
x"01fd0",-- 509
x"006e0",-- 110
x"003e0",-- 62
x"fefd0",-- -259
x"00af0",-- 175
x"00d90",-- 217
x"00b60",-- 182
x"00c50",-- 197
x"000f0",-- 15
x"ffce0",-- -50
x"febe0",-- -322
x"001e0",-- 30
x"00700",-- 112
x"ff2b0",-- -213
x"ff950",-- -107
x"ff1f0",-- -225
x"ffd80",-- -40
x"00d90",-- 217
x"ffe90",-- -23
x"002f0",-- 47
x"ff4e0",-- -178
x"ff650",-- -155
x"00280",-- 40
x"ff830",-- -125
x"00160",-- 22
x"ff800",-- -128
x"ffbf0",-- -65
x"00760",-- 118
x"00440",-- 68
x"00320",-- 50
x"ff580",-- -168
x"ffef0",-- -17
x"00b90",-- 185
x"00cf0",-- 207
x"00d90",-- 217
x"ff5d0",-- -163
x"ff600",-- -160
x"ffc20",-- -62
x"ffe40",-- -28
x"006c0",-- 108
x"00050",-- 5
x"ff8f0",-- -113
x"ffd80",-- -40
x"00aa0",-- 170
x"000c0",-- 12
x"ff4e0",-- -178
x"ffb30",-- -77
x"ff7e0",-- -130
x"003c0",-- 60
x"00820",-- 130
x"00800",-- 128
x"ffe40",-- -28
x"ff600",-- -160
x"fffb0",-- -5
x"00a00",-- 160
x"005a0",-- 90
x"ffda0",-- -38
x"00b90",-- 185
x"00710",-- 113
x"01310",-- 305
x"01360",-- 310
x"01010",-- 257
x"003a0",-- 58
x"00910",-- 145
x"009b0",-- 155
x"00be0",-- 190
x"01130",-- 275
x"ffb00",-- -80
x"00850",-- 133
x"fffe0",-- -2
x"00620",-- 98
x"00390",-- 57
x"ff860",-- -122
x"ff950",-- -107
x"fede0",-- -290
x"00370",-- 55
x"00030",-- 3
x"ffe50",-- -27
x"ff950",-- -107
x"ff7c0",-- -132
x"00280",-- 40
x"00520",-- 82
x"fff40",-- -12
x"00480",-- 72
x"00210",-- 33
x"00910",-- 145
x"00cd0",-- 205
x"00410",-- 65
x"00530",-- 83
x"00440",-- 68
x"00490",-- 73
x"fffd0",-- -3
x"00460",-- 70
x"008f0",-- 143
x"00070",-- 7
x"ffc20",-- -62
x"00020",-- 2
x"ffc10",-- -63
x"00620",-- 98
x"fff30",-- -13
x"fff80",-- -8
x"ff950",-- -107
x"ff900",-- -112
x"ffc60",-- -58
x"00530",-- 83
x"00210",-- 33
x"ffa30",-- -93
x"ffdd0",-- -35
x"ffdb0",-- -37
x"001b0",-- 27
x"00410",-- 65
x"00530",-- 83
x"00320",-- 50
x"00530",-- 83
x"00ac0",-- 172
x"01350",-- 309
x"012e0",-- 302
x"00b90",-- 185
x"00840",-- 132
x"00530",-- 83
x"00960",-- 150
x"00a30",-- 163
x"00110",-- 17
x"000c0",-- 12
x"00890",-- 137
x"00b90",-- 185
x"008e0",-- 142
x"002a0",-- 42
x"ffa60",-- -90
x"ff6f0",-- -145
x"ffe50",-- -27
x"ffd80",-- -40
x"ffb80",-- -72
x"00170",-- 23
x"ffea0",-- -22
x"00870",-- 135
x"006e0",-- 110
x"ffec0",-- -20
x"ff970",-- -105
x"ff6c0",-- -148
x"ff670",-- -153
x"ff990",-- -103
x"000f0",-- 15
x"001c0",-- 28
x"ffc10",-- -63
x"ffcc0",-- -52
x"fff60",-- -10
x"000c0",-- 12
x"ffd80",-- -40
x"ff8f0",-- -113
x"ff6a0",-- -150
x"ffdd0",-- -35
x"ffd50",-- -43
x"ffcc0",-- -52
x"fff80",-- -8
x"ff440",-- -188
x"ff8d0",-- -115
x"ff940",-- -108
x"ffd00",-- -48
x"ffe40",-- -28
x"ff950",-- -107
x"ffb50",-- -75
x"00120",-- 18
x"003e0",-- 62
x"00000",-- 0
x"00190",-- 25
x"ffdd0",-- -35
x"fffb0",-- -5
x"00140",-- 20
x"00a80",-- 168
x"00d50",-- 213
x"00960",-- 150
x"00d40",-- 212
x"01060",-- 262
x"01300",-- 304
x"00d70",-- 215
x"00ac0",-- 172
x"00530",-- 83
x"005d0",-- 93
x"008c0",-- 140
x"00660",-- 102
x"00370",-- 55
x"ff670",-- -153
x"ff950",-- -107
x"ffd80",-- -40
x"ffad0",-- -83
x"ff600",-- -160
x"ff100",-- -240
x"ff2e0",-- -210
x"ff530",-- -173
x"ff6a0",-- -150
x"ff600",-- -160
x"ff580",-- -168
x"ff070",-- -249
x"ff650",-- -155
x"ffee0",-- -18
x"00430",-- 67
x"00000",-- 0
x"ffdb0",-- -37
x"00080",-- 8
x"00750",-- 117
x"00840",-- 132
x"004e0",-- 78
x"00640",-- 100
x"000a0",-- 10
x"001e0",-- 30
x"00200",-- 32
x"003f0",-- 63
x"ffee0",-- -18
x"ffa60",-- -90
x"ff9f0",-- -97
x"ffce0",-- -50
x"ffb80",-- -72
x"ff990",-- -103
x"ff990",-- -103
x"ff990",-- -103
x"ffbd0",-- -67
x"ff850",-- -123
x"ffc20",-- -62
x"ff4e0",-- -178
x"ff650",-- -155
x"ff3a0",-- -198
x"ff790",-- -135
x"ff6c0",-- -148
x"ff450",-- -187
x"ffc60",-- -58
x"ff990",-- -103
x"ffee0",-- -18
x"ffa30",-- -93
x"00050",-- 5
x"ffce0",-- -50
x"ffd80",-- -40
x"00070",-- 7
x"00120",-- 18
x"006e0",-- 110
x"ffe20",-- -30
x"00210",-- 33
x"00140",-- 20
x"00530",-- 83
x"fff80",-- -8
x"001c0",-- 28
x"fffb0",-- -5
x"000d0",-- 13
x"00120",-- 18
x"002b0",-- 43
x"005a0",-- 90
x"000f0",-- 15
x"00500",-- 80
x"00170",-- 23
x"00570",-- 87
x"ffea0",-- -22
x"ffda0",-- -38
x"ffad0",-- -83
x"ffa80",-- -88
x"ffe90",-- -23
x"ffdf0",-- -33
x"00530",-- 83
x"ffee0",-- -18
x"003e0",-- 62
x"001e0",-- 30
x"005c0",-- 92
x"00260",-- 38
x"001c0",-- 28
x"fff30",-- -13
x"fff40",-- -12
x"003e0",-- 62
x"00300",-- 48
x"005d0",-- 93
x"00120",-- 18
x"000f0",-- 15
x"ffbd0",-- -67
x"002b0",-- 43
x"ffe00",-- -32
x"000c0",-- 12
x"ffee0",-- -18
x"fff10",-- -15
x"004b0",-- 75
x"002b0",-- 43
x"002b0",-- 43
x"ffd10",-- -47
x"fff60",-- -10
x"ff940",-- -108
x"ffe50",-- -27
x"ffa90",-- -87
x"ffe40",-- -28
x"ffd80",-- -40
x"ffd10",-- -47
x"00490",-- 73
x"00440",-- 68
x"004b0",-- 75
x"ffbf0",-- -65
x"fff10",-- -15
x"ff600",-- -160
x"ffdb0",-- -37
x"ffa30",-- -93
x"fffe0",-- -2
x"00210",-- 33
x"ffe20",-- -30
x"005c0",-- 92
x"00500",-- 80
x"003a0",-- 58
x"ffa60",-- -90
x"ffd10",-- -47
x"ff970",-- -105
x"ffec0",-- -20
x"00000",-- 0
x"00210",-- 33
x"003a0",-- 58
x"00120",-- 18
x"00410",-- 65
x"00120",-- 18
x"00340",-- 52
x"ff770",-- -137
x"ff9e0",-- -98
x"ffa90",-- -87
x"ffe70",-- -25
x"00460",-- 70
x"00340",-- 52
x"006b0",-- 107
x"00050",-- 5
x"00430",-- 67
x"fff40",-- -12
x"ffe50",-- -27
x"ff740",-- -140
x"ff9f0",-- -97
x"ffe50",-- -27
x"00030",-- 3
x"00390",-- 57
x"00210",-- 33
x"004e0",-- 78
x"fffe0",-- -2
x"fff30",-- -13
x"ffb70",-- -73
x"ff950",-- -107
x"ff3b0",-- -197
x"ff860",-- -122
x"ffd10",-- -47
x"00050",-- 5
x"002f0",-- 47
x"00160",-- 22
x"007d0",-- 125
x"00250",-- 37
x"00000",-- 0
x"ffdf0",-- -33
x"ffc90",-- -55
x"ffb50",-- -75
x"ffe40",-- -28
x"00210",-- 33
x"00530",-- 83
x"00570",-- 87
x"00410",-- 65
x"00690",-- 105
x"ffee0",-- -18
x"ffd50",-- -43
x"ff7c0",-- -132
x"ffc10",-- -63
x"ff9f0",-- -97
x"ffb80",-- -72
x"00160",-- 22
x"003c0",-- 60
x"00370",-- 55
x"ffef0",-- -17
x"00020",-- 2
x"ff810",-- -127
x"ffa10",-- -95
x"ff490",-- -183
x"ffce0",-- -50
x"ffe90",-- -23
x"00190",-- 25
x"00660",-- 102
x"00910",-- 145
x"00990",-- 153
x"000f0",-- 15
x"00370",-- 55
x"ffa90",-- -87
x"fffb0",-- -5
x"ff8d0",-- -115
x"00000",-- 0
x"fff80",-- -8
x"00490",-- 73
x"00730",-- 115
x"005f0",-- 95
x"00960",-- 150
x"ffd80",-- -40
x"001e0",-- 30
x"ff8f0",-- -113
x"fff80",-- -8
x"ffa90",-- -87
x"00020",-- 2
x"00020",-- 2
x"002b0",-- 43
x"00700",-- 112
x"004b0",-- 75
x"00750",-- 117
x"ffb00",-- -80
x"fff30",-- -13
x"ff9c0",-- -100
x"00120",-- 18
x"ffee0",-- -18
x"002d0",-- 45
x"00640",-- 100
x"007d0",-- 125
x"00bc0",-- 188
x"003e0",-- 62
x"00640",-- 100
x"ff9e0",-- -98
x"fffe0",-- -2
x"ffd50",-- -43
x"002d0",-- 45
x"00160",-- 22
x"000c0",-- 12
x"00480",-- 72
x"00300",-- 48
x"00760",-- 118
x"ffdd0",-- -35
x"00000",-- 0
x"ff950",-- -107
x"fff80",-- -8
x"fff80",-- -8
x"002b0",-- 43
x"004b0",-- 75
x"00120",-- 18
x"00410",-- 65
x"00110",-- 17
x"00480",-- 72
x"ffef0",-- -17
x"00120",-- 18
x"ffd10",-- -47
x"00160",-- 22
x"002a0",-- 42
x"00690",-- 105
x"00930",-- 147
x"00580",-- 88
x"00840",-- 132
x"003f0",-- 63
x"006c0",-- 108
x"fff10",-- -15
x"000c0",-- 12
x"ffec0",-- -20
x"00110",-- 17
x"00210",-- 33
x"00530",-- 83
x"00610",-- 97
x"00160",-- 22
x"003c0",-- 60
x"00120",-- 18
x"005c0",-- 92
x"fff80",-- -8
x"00050",-- 5
x"ffdf0",-- -33
x"00250",-- 37
x"00410",-- 65
x"00350",-- 53
x"006b0",-- 107
x"003a0",-- 58
x"00640",-- 100
x"003a0",-- 58
x"00700",-- 112
x"00320",-- 50
x"00210",-- 33
x"00190",-- 25
x"003c0",-- 60
x"00410",-- 65
x"00280",-- 40
x"00370",-- 55
x"000f0",-- 15
x"002f0",-- 47
x"fffe0",-- -2
x"00210",-- 33
x"00000",-- 0
x"ffe20",-- -30
x"00000",-- 0
x"000c0",-- 12
x"00340",-- 52
x"00000",-- 0
x"00000",-- 0
x"00030",-- 3
x"001b0",-- 27
x"00000",-- 0
x"00120",-- 18
x"00080",-- 8
x"00000",-- 0
x"002d0",-- 45
x"00320",-- 50
x"004b0",-- 75
x"00140",-- 20
x"00280",-- 40
x"00120",-- 18
x"00320",-- 50
x"000d0",-- 13
x"00140",-- 20
x"00280",-- 40
x"00120",-- 18
x"00550",-- 85
x"00260",-- 38
x"00530",-- 83
x"00070",-- 7
x"00280",-- 40
x"00020",-- 2
x"fff90",-- -7
x"00000",-- 0
x"ffd30",-- -45
x"00000",-- 0
x"fff90",-- -7
x"00300",-- 48
x"000f0",-- 15
x"00300",-- 48
x"000c0",-- 12
x"00110",-- 17
x"00020",-- 2
x"00000",-- 0
x"fffb0",-- -5
x"ffe00",-- -32
x"000d0",-- 13
x"00160",-- 22
x"00460",-- 70
x"00320",-- 50
x"00280",-- 40
x"00190",-- 25
x"00120",-- 18
x"00080",-- 8
x"fff60",-- -10
x"fffe0",-- -2
x"fff80",-- -8
x"000f0",-- 15
x"000c0",-- 12
x"00320",-- 50
x"00160",-- 22
x"00050",-- 5
x"000c0",-- 12
x"fffd0",-- -3
x"00070",-- 7
x"fffd0",-- -3
x"000d0",-- 13
x"00210",-- 33
x"002a0",-- 42
x"00370",-- 55
x"003a0",-- 58
x"00350",-- 53
x"002b0",-- 43
x"00120",-- 18
x"001b0",-- 27
x"00140",-- 20
x"00210",-- 33
x"00260",-- 38
x"002b0",-- 43
x"00350",-- 53
x"002b0",-- 43
x"00370",-- 55
x"00280",-- 40
x"00190",-- 25
x"00000",-- 0
x"fff80",-- -8
x"000f0",-- 15
x"00200",-- 32
x"00440",-- 68
x"00440",-- 68
x"00460",-- 70
x"00340",-- 52
x"00410",-- 65
x"00320",-- 50
x"000d0",-- 13
x"00050",-- 5
x"00000",-- 0
x"00170",-- 23
x"00280",-- 40
x"00390",-- 57
x"00260",-- 38
x"00440",-- 68
x"00200",-- 32
x"000d0",-- 13
x"fffb0",-- -5
x"fff30",-- -13
x"00000",-- 0
x"000c0",-- 12
x"002a0",-- 42
x"001b0",-- 27
x"003c0",-- 60
x"00210",-- 33
x"00320",-- 50
x"000f0",-- 15
x"00020",-- 2
x"00080",-- 8
x"000d0",-- 13
x"002b0",-- 43
x"00280",-- 40
x"003a0",-- 58
x"00260",-- 38
x"00370",-- 55
x"00120",-- 18
x"002d0",-- 45
x"000f0",-- 15
x"fff40",-- -12
x"fffd0",-- -3
x"00000",-- 0
x"001e0",-- 30
x"00120",-- 18
x"00230",-- 35
x"001b0",-- 27
x"00250",-- 37
x"000f0",-- 15
x"00170",-- 23
x"000a0",-- 10
x"00080",-- 8
x"00160",-- 22
x"002f0",-- 47
x"003e0",-- 62
x"00370",-- 55
x"00480",-- 72
x"001e0",-- 30
x"00210",-- 33
x"00160",-- 22
x"00160",-- 22
x"00110",-- 17
x"000c0",-- 12
x"00200",-- 32
x"002d0",-- 45
x"00390",-- 57
x"00200",-- 32
x"001e0",-- 30
x"00020",-- 2
x"000d0",-- 13
x"00020",-- 2
x"fff60",-- -10
x"fff90",-- -7
x"fff90",-- -7
x"00050",-- 5
x"fff80",-- -8
x"000d0",-- 13
x"00000",-- 0
x"fff40",-- -12
x"ffee0",-- -18
x"00000",-- 0
x"fff90",-- -7
x"ffdd0",-- -35
x"ffe70",-- -25
x"ffdf0",-- -33
x"00080",-- 8
x"000f0",-- 15
x"001c0",-- 28
x"00050",-- 5
x"fff40",-- -12
x"fff10",-- -15
x"fff10",-- -15
x"00000",-- 0
x"fff40",-- -12
x"fff40",-- -12
x"ffe50",-- -27
x"00000",-- 0
x"00020",-- 2
x"fffd0",-- -3
x"fff80",-- -8
x"ffe70",-- -25
x"ffe50",-- -27
x"ffe20",-- -30
x"fff60",-- -10
x"fffb0",-- -5
x"fff40",-- -12
x"00000",-- 0
x"00080",-- 8
x"000c0",-- 12
x"000d0",-- 13
x"00000",-- 0
x"00050",-- 5
x"00080",-- 8
x"fffe0",-- -2
x"00050",-- 5
x"fff90",-- -7
x"00050",-- 5
x"00030",-- 3
x"000c0",-- 12
x"fffe0",-- -2
x"ffec0",-- -20
x"ffe20",-- -30
x"ffdf0",-- -33
x"ffee0",-- -18
x"ffee0",-- -18
x"ffe20",-- -30
x"ffda0",-- -38
x"ffe20",-- -30
x"ffdf0",-- -33
x"ffe20",-- -30
x"ffdf0",-- -33
x"ffe20",-- -30
x"ffd30",-- -45
x"ffe00",-- -32
x"ffdf0",-- -33
x"ffd80",-- -40
x"ffe50",-- -27
x"ffec0",-- -20
x"fff80",-- -8
x"ffec0",-- -20
x"ffe70",-- -25
x"ffe90",-- -23
x"ffea0",-- -22
x"fff80",-- -8
x"ffee0",-- -18
x"ffe50",-- -27
x"ffe70",-- -25
x"ffdb0",-- -37
x"ffd80",-- -40
x"ffdf0",-- -33
x"ffee0",-- -18
x"ffe00",-- -32
x"ffd30",-- -45
x"ffc40",-- -60
x"ffce0",-- -50
x"ffd10",-- -47
x"ffd50",-- -43
x"ffd50",-- -43
x"ffd30",-- -45
x"ffd80",-- -40
x"ffe00",-- -32
x"ffdf0",-- -33
x"ffdb0",-- -37
x"ffce0",-- -50
x"ffc70",-- -57
x"ffce0",-- -50
x"ffc20",-- -62
x"ffd10",-- -47
x"ffd50",-- -43
x"ffda0",-- -38
x"ffd10",-- -47
x"ffd10",-- -47
x"ffcb0",-- -53
x"ffd10",-- -47
x"ffc70",-- -57
x"ffc60",-- -58
x"ffd60",-- -42
x"ffc10",-- -63
x"ffc60",-- -58
x"ffc70",-- -57
x"ffd50",-- -43
x"ffdf0",-- -33
x"ffda0",-- -38
x"ffd60",-- -42
x"ffc90",-- -55
x"ffc20",-- -62
x"ffbf0",-- -65
x"ffc90",-- -55
x"ffc90",-- -55
x"ffcb0",-- -53
x"ffd50",-- -43
x"ffda0",-- -38
x"ffd00",-- -48
x"ffdf0",-- -33
x"ffe40",-- -28
x"ffdb0",-- -37
x"ffec0",-- -20
x"ffdb0",-- -37
x"ffd80",-- -40
x"ffdd0",-- -35
x"ffe50",-- -27
x"ffdd0",-- -35
x"ffd80",-- -40
x"ffd60",-- -42
x"ffd60",-- -42
x"ffda0",-- -38
x"ffdb0",-- -37
x"ffdb0",-- -37
x"ffdf0",-- -33
x"ffe20",-- -30
x"ffe50",-- -27
x"ffe50",-- -27
x"ffd80",-- -40
x"ffea0",-- -22
x"ffe20",-- -30
x"ffe00",-- -32
x"ffd50",-- -43
x"ffdb0",-- -37
x"ffe20",-- -30
x"ffdf0",-- -33
x"ffec0",-- -20
x"ffef0",-- -17
x"fff80",-- -8
x"ffec0",-- -20
x"ffee0",-- -18
x"ffea0",-- -22
x"ffe20",-- -30
x"fff10",-- -15
x"ffee0",-- -18
x"ffee0",-- -18
x"fffb0",-- -5
x"ffea0",-- -22
x"ffea0",-- -22
x"ffea0",-- -22
x"ffe00",-- -32
x"ffdb0",-- -37
x"ffdb0",-- -37
x"ffe40",-- -28
x"ffe50",-- -27
x"ffea0",-- -22
x"fff40",-- -12
x"ffee0",-- -18
x"ffea0",-- -22
x"ffe50",-- -27
x"ffea0",-- -22
x"ffee0",-- -18
x"ffea0",-- -22
x"ffea0",-- -22
x"ffef0",-- -17
x"fff40",-- -12
x"ffee0",-- -18
x"fffe0",-- -2
x"00000",-- 0
x"fff30",-- -13
x"fff60",-- -10
x"00000",-- 0
x"fffe0",-- -2
x"fff60",-- -10
x"fff90",-- -7
x"fffb0",-- -5
x"fffd0",-- -3
x"fffe0",-- -2
x"00000",-- 0
x"000d0",-- 13
x"00000",-- 0
x"00000",-- 0
x"00080",-- 8
x"00050",-- 5
x"00120",-- 18
x"00140",-- 20
x"00050",-- 5
x"00020",-- 2
x"00050",-- 5
x"00030",-- 3
x"00050",-- 5
x"00070",-- 7
x"000c0",-- 12
x"00030",-- 3
x"00020",-- 2
x"000c0",-- 12
x"000c0",-- 12
x"00110",-- 17
x"000c0",-- 12
x"00160",-- 22
x"001b0",-- 27
x"00170",-- 23
x"00160",-- 22
x"00120",-- 18
x"000f0",-- 15
x"00080",-- 8
x"00160",-- 22
x"00140",-- 20
x"000c0",-- 12
x"000c0",-- 12
x"00050",-- 5
x"000f0",-- 15
x"001e0",-- 30
x"00160",-- 22
x"00120",-- 18
x"000c0",-- 12
x"000c0",-- 12
x"000c0",-- 12
x"00160",-- 22
x"000f0",-- 15
x"00030",-- 3
x"00080",-- 8
x"00080",-- 8
x"001c0",-- 28
x"00140",-- 20
x"00120",-- 18
x"000d0",-- 13
x"00120",-- 18
x"000f0",-- 15
x"00000",-- 0
x"000c0",-- 12
x"00050",-- 5
x"000d0",-- 13
x"001e0",-- 30
x"001b0",-- 27
x"00120",-- 18
x"000f0",-- 15
x"00070",-- 7
x"00120",-- 18
x"000c0",-- 12
x"00070",-- 7
x"00120",-- 18
x"00020",-- 2
x"00110",-- 17
x"00120",-- 18
x"00110",-- 17
x"00080",-- 8
x"000f0",-- 15
x"00110",-- 17
x"000c0",-- 12
x"00160",-- 22
x"001b0",-- 27
x"00170",-- 23
x"000f0",-- 15
x"000a0",-- 10
x"00050",-- 5
x"00110",-- 17
x"000d0",-- 13
x"00000",-- 0
x"000a0",-- 10
x"00070",-- 7
x"000c0",-- 12
x"00110",-- 17
x"00050",-- 5
x"000c0",-- 12
x"000d0",-- 13
x"00120",-- 18
x"000c0",-- 12
x"00020",-- 2
x"00080",-- 8
x"00030",-- 3
x"00000",-- 0
x"00000",-- 0
x"00020",-- 2
x"000c0",-- 12
x"00080",-- 8
x"00050",-- 5
x"00000",-- 0
x"00020",-- 2
x"000c0",-- 12
x"000c0",-- 12
x"001b0",-- 27
x"000f0",-- 15
x"000a0",-- 10
x"000a0",-- 10
x"00050",-- 5
x"000f0",-- 15
x"00070",-- 7
x"00140",-- 20
x"00160",-- 22
x"00050",-- 5
x"00070",-- 7
x"00030",-- 3
x"00080",-- 8
x"00030",-- 3
x"00000",-- 0
x"00080",-- 8
x"00000",-- 0
x"00020",-- 2
x"00080",-- 8
x"00000",-- 0
x"00000",-- 0
x"00050",-- 5
x"00050",-- 5
x"00020",-- 2
x"00070",-- 7
x"00030",-- 3
x"00020",-- 2
x"00020",-- 2
x"00080",-- 8
x"000f0",-- 15
x"00110",-- 17
x"000c0",-- 12
x"00080",-- 8
x"000d0",-- 13
x"00070",-- 7
x"000c0",-- 12
x"00070",-- 7
x"00110",-- 17
x"00160",-- 22
x"00120",-- 18
x"00120",-- 18
x"00160",-- 22
x"000f0",-- 15
x"00030",-- 3
x"000f0",-- 15
x"00120",-- 18
x"00140",-- 20
x"001c0",-- 28
x"00280",-- 40
x"00200",-- 32
x"00210",-- 33
x"001b0",-- 27
x"000a0",-- 10
x"00190",-- 25
x"00160",-- 22
x"00170",-- 23
x"00160",-- 22
x"00110",-- 17
x"00080",-- 8
x"000c0",-- 12
x"00070",-- 7
x"000f0",-- 15
x"00140",-- 20
x"00070",-- 7
x"000c0",-- 12
x"00050",-- 5
x"00050",-- 5
x"00050",-- 5
x"00050",-- 5
x"000c0",-- 12
x"00050",-- 5
x"000d0",-- 13
x"000f0",-- 15
x"00110",-- 17
x"00140",-- 20
x"00190",-- 25
x"00160",-- 22
x"000c0",-- 12
x"000a0",-- 10
x"00120",-- 18
x"00190",-- 25
x"00210",-- 33
x"001e0",-- 30
x"001b0",-- 27
x"001c0",-- 28
x"001c0",-- 28
x"002b0",-- 43
x"000f0",-- 15
x"00250",-- 37
x"001c0",-- 28
x"00260",-- 38
x"00280",-- 40
x"001e0",-- 30
x"00370",-- 55
x"00210",-- 33
x"00320",-- 50
x"002f0",-- 47
x"002a0",-- 42
x"003e0",-- 62
x"00430",-- 67
x"00350",-- 53
x"00320",-- 50
x"002d0",-- 45
x"002f0",-- 47
x"00370",-- 55
x"00350",-- 53
x"00370",-- 55
x"00210",-- 33
x"00210",-- 33
x"00280",-- 40
x"00250",-- 37
x"001c0",-- 28
x"00120",-- 18
x"00140",-- 20
x"001e0",-- 30
x"001b0",-- 27
x"00170",-- 23
x"00260",-- 38
x"00190",-- 25
x"00280",-- 40
x"00280",-- 40
x"00280",-- 40
x"002b0",-- 43
x"00250",-- 37
x"00210",-- 33
x"00280",-- 40
x"00250",-- 37
x"00230",-- 35
x"002f0",-- 47
x"00210",-- 33
x"001b0",-- 27
x"00210",-- 33
x"002d0",-- 45
x"00280",-- 40
x"00200",-- 32
x"00170",-- 23
x"000f0",-- 15
x"000f0",-- 15
x"000d0",-- 13
x"001c0",-- 28
x"001b0",-- 27
x"001b0",-- 27
x"001b0",-- 27
x"000d0",-- 13
x"00110",-- 17
x"001b0",-- 27
x"00120",-- 18
x"000c0",-- 12
x"000c0",-- 12
x"00120",-- 18
x"00160",-- 22
x"000d0",-- 13
x"000f0",-- 15
x"00170",-- 23
x"000f0",-- 15
x"001e0",-- 30
x"000d0",-- 13
x"00000",-- 0
x"000c0",-- 12
x"00050",-- 5
x"00050",-- 5
x"000c0",-- 12
x"00050",-- 5
x"00190",-- 25
x"001b0",-- 27
x"00000",-- 0
x"00080",-- 8
x"00030",-- 3
x"00000",-- 0
x"00020",-- 2
x"00000",-- 0
x"00020",-- 2
x"00000",-- 0
x"00080",-- 8
x"00030",-- 3
x"00110",-- 17
x"000f0",-- 15
x"00000",-- 0
x"00070",-- 7
x"00000",-- 0
x"00020",-- 2
x"00110",-- 17
x"00020",-- 2
x"00080",-- 8
x"00120",-- 18
x"00070",-- 7
x"00070",-- 7
x"00020",-- 2
x"fffe0",-- -2
x"00000",-- 0
x"00000",-- 0
x"fff40",-- -12
x"fff80",-- -8
x"fff10",-- -15
x"fff80",-- -8
x"00000",-- 0
x"fffb0",-- -5
x"fffe0",-- -2
x"fff30",-- -13
x"fff60",-- -10
x"fff40",-- -12
x"ffee0",-- -18
x"fffe0",-- -2
x"fffb0",-- -5
x"ffef0",-- -17
x"fff10",-- -15
x"ffe50",-- -27
x"fff40",-- -12
x"fffb0",-- -5
x"fff80",-- -8
x"fff40",-- -12
x"fff30",-- -13
x"ffee0",-- -18
x"fff80",-- -8
x"fffb0",-- -5
x"fffe0",-- -2
x"fffd0",-- -3
x"fff30",-- -13
x"00000",-- 0
x"fffb0",-- -5
x"fff60",-- -10
x"fff10",-- -15
x"fffd0",-- -3
x"00030",-- 3
x"00030",-- 3
x"00080",-- 8
x"fffe0",-- -2
x"ffee0",-- -18
x"00000",-- 0
x"fffe0",-- -2
x"fff10",-- -15
x"fff40",-- -12
x"ffee0",-- -18
x"fff60",-- -10
x"ffec0",-- -20
x"ffee0",-- -18
x"ffee0",-- -18
x"ffea0",-- -22
x"ffdf0",-- -33
x"ffe00",-- -32
x"ffe70",-- -25
x"ffe50",-- -27
x"ffee0",-- -18
x"fff30",-- -13
x"fff80",-- -8
x"fff90",-- -7
x"00000",-- 0
x"ffe50",-- -27
x"00000",-- 0
x"fff10",-- -15
x"fffe0",-- -2
x"ffec0",-- -20
x"ffe20",-- -30
x"fff80",-- -8
x"ffe50",-- -27
x"fffb0",-- -5
x"ffee0",-- -18
x"ffe90",-- -23
x"ffe20",-- -30
x"ffee0",-- -18
x"ffdf0",-- -33
x"fffe0",-- -2
x"fffe0",-- -2
x"ffdd0",-- -35
x"fff40",-- -12
x"fff40",-- -12
x"00000",-- 0
x"fff80",-- -8
x"fffb0",-- -5
x"ffee0",-- -18
x"fff10",-- -15
x"00000",-- 0
x"fff90",-- -7
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fffe0",-- -2
x"00020",-- 2
x"00000",-- 0
x"fff60",-- -10
x"fff40",-- -12
x"fff60",-- -10
x"ffea0",-- -22
x"ffef0",-- -17
x"ffea0",-- -22
x"ffee0",-- -18
x"fffb0",-- -5
x"00050",-- 5
x"fffd0",-- -3
x"fffb0",-- -5
x"00000",-- 0
x"fff40",-- -12
x"00000",-- 0
x"fff10",-- -15
x"fff40",-- -12
x"00020",-- 2
x"fffd0",-- -3
x"fff90",-- -7
x"fffd0",-- -3
x"00000",-- 0
x"fff80",-- -8
x"fffb0",-- -5
x"fffe0",-- -2
x"fffe0",-- -2
x"00020",-- 2
x"00000",-- 0
x"00000",-- 0
x"00020",-- 2
x"00020",-- 2
x"00000",-- 0
x"fff90",-- -7
x"fffe0",-- -2
x"fff80",-- -8
x"00000",-- 0
x"00020",-- 2
x"00000",-- 0
x"fffd0",-- -3
x"00000",-- 0
x"00000",-- 0
x"fffd0",-- -3
x"fffb0",-- -5
x"fff40",-- -12
x"fffb0",-- -5
x"00000",-- 0
x"00050",-- 5
x"fffe0",-- -2
x"fffe0",-- -2
x"ffee0",-- -18
x"fffe0",-- -2
x"fff80",-- -8
x"ffef0",-- -17
x"ffea0",-- -22
x"ffe40",-- -28
x"ffe90",-- -23
x"fff10",-- -15
x"fff40",-- -12
x"ffe50",-- -27
x"fff10",-- -15
x"ffea0",-- -22
x"ffe90",-- -23
x"ffdd0",-- -35
x"ffe20",-- -30
x"ffdf0",-- -33
x"ffe20",-- -30
x"ffdf0",-- -33
x"ffe20",-- -30
x"ffee0",-- -18
x"ffe90",-- -23
x"ffdd0",-- -35
x"ffdb0",-- -37
x"ffe40",-- -28
x"ffe20",-- -30
x"ffe50",-- -27
x"ffee0",-- -18
x"ffdd0",-- -35
x"ffdd0",-- -35
x"ffe70",-- -25
x"ffe50",-- -27
x"ffee0",-- -18
x"fff10",-- -15
x"fff40",-- -12
x"fff60",-- -10
x"fff60",-- -10
x"ffea0",-- -22
x"ffe40",-- -28
x"ffea0",-- -22
x"ffe20",-- -30
x"ffee0",-- -18
x"ffe50",-- -27
x"ffe20",-- -30
x"ffe50",-- -27
x"ffe20",-- -30
x"ffd60",-- -42
x"ffd10",-- -47
x"ffea0",-- -22
x"ffe20",-- -30
x"ffea0",-- -22
x"fff10",-- -15
x"ffea0",-- -22
x"ffe70",-- -25
x"ffef0",-- -17
x"ffee0",-- -18
x"ffe90",-- -23
x"ffe20",-- -30
x"ffea0",-- -22
x"ffee0",-- -18
x"ffe20",-- -30
x"ffea0",-- -22
x"ffec0",-- -20
x"fff10",-- -15
x"fff90",-- -7
x"ffea0",-- -22
x"ffe50",-- -27
x"ffd80",-- -40
x"ffd50",-- -43
x"ffdf0",-- -33
x"ffdb0",-- -37
x"ffe40",-- -28
x"ffdf0",-- -33
x"ffea0",-- -22
x"ffe20",-- -30
x"ffdd0",-- -35
x"ffdf0",-- -33
x"fff10",-- -15
x"ffea0",-- -22
x"ffe00",-- -32
x"ffe20",-- -30
x"fff10",-- -15
x"fff30",-- -13
x"ffe90",-- -23
x"ffea0",-- -22
x"ffe20",-- -30
x"ffe50",-- -27
x"ffef0",-- -17
x"ffec0",-- -20
x"ffee0",-- -18
x"ffe20",-- -30
x"ffee0",-- -18
x"ffee0",-- -18
x"ffdb0",-- -37
x"ffee0",-- -18
x"ffea0",-- -22
x"ffe40",-- -28
x"ffee0",-- -18
x"ffee0",-- -18
x"fff10",-- -15
x"fff40",-- -12
x"ffe50",-- -27
x"ffec0",-- -20
x"fff80",-- -8
x"fff90",-- -7
x"00000",-- 0
x"fff80",-- -8
x"fffe0",-- -2
x"fffe0",-- -2
x"fff80",-- -8
x"fffe0",-- -2
x"00000",-- 0
x"fff40",-- -12
x"00000",-- 0
x"fffe0",-- -2
x"fffe0",-- -2
x"00020",-- 2
x"00020",-- 2
x"00020",-- 2
x"00020",-- 2
x"000f0",-- 15
x"00110",-- 17
x"00120",-- 18
x"001c0",-- 28
x"00140",-- 20
x"00190",-- 25
x"00110",-- 17
x"000c0",-- 12
x"00080",-- 8
x"000c0",-- 12
x"00110",-- 17
x"000f0",-- 15
x"00120",-- 18
x"00020",-- 2
x"00000",-- 0
x"00020",-- 2
x"00030",-- 3
x"00080",-- 8
x"00080",-- 8
x"000c0",-- 12
x"00080",-- 8
x"fffe0",-- -2
x"00000",-- 0
x"00020",-- 2
x"00050",-- 5
x"00050",-- 5
x"00080",-- 8
x"00070",-- 7
x"00000",-- 0
x"00000",-- 0
x"fffe0",-- -2
x"fff40",-- -12
x"fff10",-- -15
x"ffe50",-- -27
x"ffee0",-- -18
x"fff40",-- -12
x"00000",-- 0
x"fff40",-- -12
x"00000",-- 0
x"fff40",-- -12
x"000f0",-- 15
x"00070",-- 7
x"fff40",-- -12
x"fff80",-- -8
x"ffc20",-- -62
x"00000",-- 0
x"00a00",-- 160
x"01bd0",-- 445
x"018a0",-- 394
x"ff2b0",-- -213
x"fd270",-- -729
x"fe570",-- -425
x"00c80",-- 200
x"017b0",-- 379
x"00b20",-- 178
x"ff810",-- -127
x"fee90",-- -279
x"00af0",-- 175
x"02b40",-- 692
x"013a0",-- 314
x"fdf90",-- -519
x"fc7a0",-- -902
x"fe020",-- -510
x"00b10",-- 177
x"02570",-- 599
x"01c70",-- 455
x"00350",-- 53
x"ffe50",-- -27
x"00eb0",-- 235
x"015e0",-- 350
x"00890",-- 137
x"ff170",-- -233
x"fddf0",-- -545
x"febc0",-- -324
x"00c50",-- 197
x"01b50",-- 437
x"010e0",-- 270
x"003a0",-- 58
x"00070",-- 7
x"003e0",-- 62
x"00230",-- 35
x"ff790",-- -135
x"feac0",-- -340
x"febe0",-- -322
x"ffce0",-- -50
x"00b40",-- 180
x"01290",-- 297
x"00f40",-- 244
x"006c0",-- 108
x"00410",-- 65
x"00700",-- 112
x"00480",-- 72
x"ff920",-- -110
x"ff1f0",-- -225
x"ff600",-- -160
x"00230",-- 35
x"00d50",-- 213
x"00f90",-- 249
x"00910",-- 145
x"00210",-- 33
x"fffb0",-- -5
x"ffe90",-- -23
x"ffb50",-- -75
x"ff6d0",-- -147
x"ff450",-- -187
x"ff8a0",-- -118
x"00370",-- 55
x"00cf0",-- 207
x"00e80",-- 232
x"009d0",-- 157
x"005f0",-- 95
x"002d0",-- 45
x"00020",-- 2
x"ffd00",-- -48
x"ff9c0",-- -100
x"ffab0",-- -85
x"fff10",-- -15
x"00610",-- 97
x"00a80",-- 168
x"00940",-- 148
x"00550",-- 85
x"00200",-- 32
x"ffe50",-- -27
x"ffbc0",-- -68
x"ff830",-- -125
x"ff710",-- -143
x"ffbc0",-- -68
x"002f0",-- 47
x"008f0",-- 143
x"00ac0",-- 172
x"00960",-- 150
x"00700",-- 112
x"004d0",-- 77
x"00160",-- 22
x"ffea0",-- -22
x"ffc90",-- -55
x"ffbf0",-- -65
x"000a0",-- 10
x"006b0",-- 107
x"007a0",-- 122
x"00700",-- 112
x"00440",-- 68
x"00230",-- 35
x"00080",-- 8
x"ffe20",-- -30
x"ffb50",-- -75
x"ff9c0",-- -100
x"ffc20",-- -62
x"000d0",-- 13
x"00550",-- 85
x"00760",-- 118
x"007b0",-- 123
x"00570",-- 87
x"00370",-- 55
x"00210",-- 33
x"fffd0",-- -3
x"ffcc0",-- -52
x"ffc60",-- -58
x"ffe50",-- -27
x"00230",-- 35
x"005c0",-- 92
x"00660",-- 102
x"00440",-- 68
x"000f0",-- 15
x"00000",-- 0
x"ffdf0",-- -33
x"ffd50",-- -43
x"ffb50",-- -75
x"ffb30",-- -77
x"ffe50",-- -27
x"001b0",-- 27
x"00640",-- 100
x"00660",-- 102
x"00300",-- 48
x"00050",-- 5
x"fff10",-- -15
x"ffe00",-- -32
x"ffdb0",-- -37
x"ffda0",-- -38
x"ffd60",-- -42
x"ffee0",-- -18
x"001e0",-- 30
x"00320",-- 50
x"003e0",-- 62
x"001b0",-- 27
x"ffe20",-- -30
x"ffc20",-- -62
x"ffc20",-- -62
x"ffce0",-- -50
x"ffe50",-- -27
x"00050",-- 5
x"00140",-- 20
x"003c0",-- 60
x"003e0",-- 62
x"004b0",-- 75
x"00370",-- 55
x"00000",-- 0
x"fff40",-- -12
x"ffee0",-- -18
x"00000",-- 0
x"00210",-- 33
x"00340",-- 52
x"00280",-- 40
x"00190",-- 25
x"000d0",-- 13
x"00160",-- 22
x"00210",-- 33
x"00080",-- 8
x"ffef0",-- -17
x"ffdd0",-- -35
x"fff10",-- -15
x"001e0",-- 30
x"003a0",-- 58
x"003a0",-- 58
x"00320",-- 50
x"00260",-- 38
x"00260",-- 38
x"00410",-- 65
x"00250",-- 37
x"000f0",-- 15
x"00050",-- 5
x"00080",-- 8
x"001c0",-- 28
x"003f0",-- 63
x"00440",-- 68
x"00200",-- 32
x"00190",-- 25
x"000f0",-- 15
x"00120",-- 18
x"00120",-- 18
x"fffb0",-- -5
x"fff10",-- -15
x"fff40",-- -12
x"00020",-- 2
x"002b0",-- 43
x"002d0",-- 45
x"002d0",-- 45
x"00200",-- 32
x"00120",-- 18
x"001c0",-- 28
x"00110",-- 17
x"00020",-- 2
x"ffec0",-- -20
x"fffe0",-- -2
x"000d0",-- 13
x"00170",-- 23
x"00200",-- 32
x"00120",-- 18
x"00080",-- 8
x"fff80",-- -8
x"fffb0",-- -5
x"fff80",-- -8
x"ffee0",-- -18
x"fffe0",-- -2
x"00000",-- 0
x"00110",-- 17
x"00250",-- 37
x"001c0",-- 28
x"000f0",-- 15
x"00080",-- 8
x"fffe0",-- -2
x"fff60",-- -10
x"ffee0",-- -18
x"ffdd0",-- -35
x"fff40",-- -12
x"fff60",-- -10
x"fff40",-- -12
x"00020",-- 2
x"fffd0",-- -3
x"fff60",-- -10
x"fff10",-- -15
x"ffee0",-- -18
x"ffe50",-- -27
x"fff80",-- -8
x"fffe0",-- -2
x"fff90",-- -7
x"000a0",-- 10
x"000f0",-- 15
x"00140",-- 20
x"00210",-- 33
x"00190",-- 25
x"000a0",-- 10
x"00080",-- 8
x"00020",-- 2
x"00000",-- 0
x"fffe0",-- -2
x"00000",-- 0
x"00160",-- 22
x"00120",-- 18
x"00190",-- 25
x"00050",-- 5
x"fffb0",-- -5
x"00020",-- 2
x"00030",-- 3
x"00050",-- 5
x"00080",-- 8
x"00070",-- 7
x"000f0",-- 15
x"00190",-- 25
x"00160",-- 22
x"001e0",-- 30
x"00140",-- 20
x"00050",-- 5
x"fff90",-- -7
x"00000",-- 0
x"00050",-- 5
x"fff60",-- -10
x"ffea0",-- -22
x"fff10",-- -15
x"fff40",-- -12
x"00000",-- 0
x"00000",-- 0
x"ffec0",-- -20
x"ffe40",-- -28
x"ffd30",-- -45
x"ffda0",-- -38
x"ffe50",-- -27
x"fff10",-- -15
x"ffee0",-- -18
x"ffef0",-- -17
x"00030",-- 3
x"00000",-- 0
x"fffb0",-- -5
x"ffe40",-- -28
x"ffc90",-- -55
x"ffc90",-- -55
x"ffdd0",-- -35
x"fff10",-- -15
x"ffdf0",-- -33
x"ffdf0",-- -33
x"ffd80",-- -40
x"ffdf0",-- -33
x"ffe50",-- -27
x"ffd80",-- -40
x"ffdb0",-- -37
x"ffd80",-- -40
x"ffd30",-- -45
x"ffdd0",-- -35
x"ffee0",-- -18
x"fff10",-- -15
x"fff30",-- -13
x"fff30",-- -13
x"fffb0",-- -5
x"00000",-- 0
x"fffe0",-- -2
x"ffee0",-- -18
x"ffe40",-- -28
x"ffec0",-- -20
x"ffef0",-- -17
x"ffee0",-- -18
x"ffe70",-- -25
x"fff90",-- -7
x"fffd0",-- -3
x"fff80",-- -8
x"fffe0",-- -2
x"ffef0",-- -17
x"fffb0",-- -5
x"fff90",-- -7
x"ffec0",-- -20
x"fff10",-- -15
x"fff40",-- -12
x"ffec0",-- -20
x"fff60",-- -10
x"fff10",-- -15
x"ffef0",-- -17
x"fff80",-- -8
x"ffe50",-- -27
x"ffdf0",-- -33
x"ffe20",-- -30
x"ffe40",-- -28
x"ffe20",-- -30
x"ffd50",-- -43
x"ffd80",-- -40
x"ffe50",-- -27
x"ffec0",-- -20
x"fff10",-- -15
x"ffe70",-- -25
x"ffe70",-- -25
x"ffdf0",-- -33
x"fff40",-- -12
x"00000",-- 0
x"ffee0",-- -18
x"ffea0",-- -22
x"fff60",-- -10
x"00070",-- 7
x"00000",-- 0
x"ffea0",-- -22
x"ffea0",-- -22
x"ffe50",-- -27
x"ffee0",-- -18
x"ffe90",-- -23
x"ffe50",-- -27
x"fff10",-- -15
x"ffef0",-- -17
x"ffe70",-- -25
x"ffe50",-- -27
x"ffef0",-- -17
x"ffea0",-- -22
x"ffea0",-- -22
x"ffe50",-- -27
x"ffdf0",-- -33
x"ffea0",-- -22
x"fff40",-- -12
x"ffef0",-- -17
x"fff40",-- -12
x"ffea0",-- -22
x"ffef0",-- -17
x"fffe0",-- -2
x"ffe90",-- -23
x"ffee0",-- -18
x"ffe90",-- -23
x"ffee0",-- -18
x"fff30",-- -13
x"fff60",-- -10
x"fffb0",-- -5
x"fff10",-- -15
x"ffef0",-- -17
x"fff90",-- -7
x"fff10",-- -15
x"ffe90",-- -23
x"ffee0",-- -18
x"ffdd0",-- -35
x"ffdb0",-- -37
x"ffe20",-- -30
x"ffdd0",-- -35
x"ffd50",-- -43
x"ffdf0",-- -33
x"ffea0",-- -22
x"ffe90",-- -23
x"ffe70",-- -25
x"ffdd0",-- -35
x"ffe00",-- -32
x"ffdb0",-- -37
x"ffe50",-- -27
x"ffea0",-- -22
x"ffe70",-- -25
x"ffdd0",-- -35
x"ffdd0",-- -35
x"ffda0",-- -38
x"ffea0",-- -22
x"ffdb0",-- -37
x"ffcc0",-- -52
x"ffd80",-- -40
x"ffe20",-- -30
x"ffee0",-- -18
x"ffe50",-- -27
x"ffe20",-- -30
x"ffd80",-- -40
x"ffe20",-- -30
x"ffe70",-- -25
x"ffe90",-- -23
x"ffdf0",-- -33
x"ffdb0",-- -37
x"ffdf0",-- -33
x"ffe50",-- -27
x"ffdb0",-- -37
x"ffda0",-- -38
x"ffdd0",-- -35
x"ffd60",-- -42
x"ffdb0",-- -37
x"ffdd0",-- -35
x"ffe00",-- -32
x"ffdf0",-- -33
x"ffe20",-- -30
x"ffdf0",-- -33
x"ffda0",-- -38
x"ffd50",-- -43
x"ffd80",-- -40
x"ffe00",-- -32
x"ffda0",-- -38
x"ffd50",-- -43
x"ffce0",-- -50
x"ffd10",-- -47
x"ffd80",-- -40
x"ffd10",-- -47
x"ffc90",-- -55
x"ffd30",-- -45
x"ffe20",-- -30
x"ffdf0",-- -33
x"ffd60",-- -42
x"ffdb0",-- -37
x"ffd50",-- -43
x"ffe50",-- -27
x"ffee0",-- -18
x"ffdf0",-- -33
x"ffea0",-- -22
x"ffea0",-- -22
x"ffe90",-- -23
x"ffee0",-- -18
x"ffe50",-- -27
x"ffea0",-- -22
x"ffe90",-- -23
x"fffb0",-- -5
x"fffb0",-- -5
x"00000",-- 0
x"00070",-- 7
x"fff90",-- -7
x"00020",-- 2
x"fffd0",-- -3
x"fff90",-- -7
x"00030",-- 3
x"fffd0",-- -3
x"00020",-- 2
x"00050",-- 5
x"fff40",-- -12
x"fffd0",-- -3
x"00000",-- 0
x"00000",-- 0
x"00020",-- 2
x"00000",-- 0
x"fff40",-- -12
x"fff10",-- -15
x"fff90",-- -7
x"00020",-- 2
x"fffb0",-- -5
x"fff60",-- -10
x"fff10",-- -15
x"fffd0",-- -3
x"00020",-- 2
x"fffe0",-- -2
x"fffe0",-- -2
x"fffb0",-- -5
x"00000",-- 0
x"fffe0",-- -2
x"fffb0",-- -5
x"fff80",-- -8
x"fff80",-- -8
x"00080",-- 8
x"00080",-- 8
x"00080",-- 8
x"00020",-- 2
x"00020",-- 2
x"00050",-- 5
x"00020",-- 2
x"00030",-- 3
x"00020",-- 2
x"00000",-- 0
x"fffe0",-- -2
x"00020",-- 2
x"00020",-- 2
x"00030",-- 3
x"00020",-- 2
x"00050",-- 5
x"000f0",-- 15
x"00080",-- 8
x"00140",-- 20
x"001b0",-- 27
x"00170",-- 23
x"001b0",-- 27
x"00140",-- 20
x"001b0",-- 27
x"001b0",-- 27
x"00110",-- 17
x"00080",-- 8
x"00170",-- 23
x"00170",-- 23
x"00160",-- 22
x"001e0",-- 30
x"00160",-- 22
x"00120",-- 18
x"001b0",-- 27
x"00170",-- 23
x"000f0",-- 15
x"00140",-- 20
x"00160",-- 22
x"00080",-- 8
x"000d0",-- 13
x"00120",-- 18
x"00120",-- 18
x"000f0",-- 15
x"000f0",-- 15
x"00160",-- 22
x"00170",-- 23
x"001c0",-- 28
x"00120",-- 18
x"000f0",-- 15
x"00020",-- 2
x"000a0",-- 10
x"000f0",-- 15
x"00190",-- 25
x"000d0",-- 13
x"00170",-- 23
x"00280",-- 40
x"00160",-- 22
x"001b0",-- 27
x"00120",-- 18
x"000f0",-- 15
x"00170",-- 23
x"00080",-- 8
x"00080",-- 8
x"000f0",-- 15
x"000a0",-- 10
x"000f0",-- 15
x"000f0",-- 15
x"000a0",-- 10
x"00080",-- 8
x"00080",-- 8
x"00110",-- 17
x"000c0",-- 12
x"00080",-- 8
x"000c0",-- 12
x"000d0",-- 13
x"00140",-- 20
x"000c0",-- 12
x"00140",-- 20
x"00160",-- 22
x"00170",-- 23
x"00110",-- 17
x"00020",-- 2
x"00080",-- 8
x"000f0",-- 15
x"00020",-- 2
x"000c0",-- 12
x"00080",-- 8
x"fffe0",-- -2
x"000a0",-- 10
x"00050",-- 5
x"00020",-- 2
x"00020",-- 2
x"00070",-- 7
x"fffe0",-- -2
x"00070",-- 7
x"00020",-- 2
x"00000",-- 0
x"000d0",-- 13
x"00000",-- 0
x"00000",-- 0
x"00020",-- 2
x"00020",-- 2
x"00020",-- 2
x"000c0",-- 12
x"00050",-- 5
x"00020",-- 2
x"000c0",-- 12
x"000c0",-- 12
x"00000",-- 0
x"fffe0",-- -2
x"00080",-- 8
x"000a0",-- 10
x"00000",-- 0
x"fffe0",-- -2
x"00030",-- 3
x"000a0",-- 10
x"00120",-- 18
x"000f0",-- 15
x"00080",-- 8
x"00020",-- 2
x"00020",-- 2
x"00050",-- 5
x"00000",-- 0
x"fffb0",-- -5
x"00000",-- 0
x"00050",-- 5
x"000c0",-- 12
x"000d0",-- 13
x"000f0",-- 15
x"00170",-- 23
x"00210",-- 33
x"00140",-- 20
x"001b0",-- 27
x"001c0",-- 28
x"00140",-- 20
x"00200",-- 32
x"001b0",-- 27
x"00250",-- 37
x"00210",-- 33
x"00210",-- 33
x"00210",-- 33
x"00230",-- 35
x"002b0",-- 43
x"00280",-- 40
x"00210",-- 33
x"00170",-- 23
x"001e0",-- 30
x"001b0",-- 27
x"00250",-- 37
x"002b0",-- 43
x"00250",-- 37
x"00280",-- 40
x"002a0",-- 42
x"00260",-- 38
x"00230",-- 35
x"00280",-- 40
x"00370",-- 55
x"00340",-- 52
x"00280",-- 40
x"00280",-- 40
x"00280",-- 40
x"002b0",-- 43
x"00200",-- 32
x"00250",-- 37
x"002d0",-- 45
x"002f0",-- 47
x"002f0",-- 47
x"00210",-- 33
x"00280",-- 40
x"00230",-- 35
x"00280",-- 40
x"00280",-- 40
x"00260",-- 38
x"00260",-- 38
x"00210",-- 33
x"00140",-- 20
x"001e0",-- 30
x"001e0",-- 30
x"00120",-- 18
x"00210",-- 33
x"00250",-- 37
x"002f0",-- 47
x"002a0",-- 42
x"002f0",-- 47
x"00230",-- 35
x"00210",-- 33
x"002a0",-- 42
x"00250",-- 37
x"00260",-- 38
x"00210",-- 33
x"00300",-- 48
x"00280",-- 40
x"00250",-- 37
x"001e0",-- 30
x"001e0",-- 30
x"002d0",-- 45
x"002b0",-- 43
x"00200",-- 32
x"00120",-- 18
x"00110",-- 17
x"00080",-- 8
x"00080",-- 8
x"fffe0",-- -2
x"00030",-- 3
x"00020",-- 2
x"00000",-- 0
x"00000",-- 0
x"fff80",-- -8
x"fff80",-- -8
x"00000",-- 0
x"00000",-- 0
x"fffe0",-- -2
x"00000",-- 0
x"fffb0",-- -5
x"00000",-- 0
x"00020",-- 2
x"00050",-- 5
x"00030",-- 3
x"00020",-- 2
x"00000",-- 0
x"fff80",-- -8
x"fffd0",-- -3
x"00000",-- 0
x"000a0",-- 10
x"000c0",-- 12
x"00000",-- 0
x"00000",-- 0
x"00000",-- 0
x"fffe0",-- -2
x"00000",-- 0
x"00050",-- 5
x"00000",-- 0
x"fffb0",-- -5
x"00000",-- 0
x"fffe0",-- -2
x"00000",-- 0
x"fffd0",-- -3
x"00050",-- 5
x"00080",-- 8
x"00020",-- 2
x"fffb0",-- -5
x"fff80",-- -8
x"00000",-- 0
x"fffe0",-- -2
x"00000",-- 0
x"00020",-- 2
x"00000",-- 0
x"fffe0",-- -2
x"fff90",-- -7
x"fffe0",-- -2
x"fff80",-- -8
x"00000",-- 0
x"00080",-- 8
x"000c0",-- 12
x"00080",-- 8
x"00000",-- 0
x"fff80",-- -8
x"00000",-- 0
x"00000",-- 0
x"00030",-- 3
x"00050",-- 5
x"00020",-- 2
x"fffb0",-- -5
x"fff40",-- -12
x"fffe0",-- -2
x"fffd0",-- -3
x"fffe0",-- -2
x"fff60",-- -10
x"00000",-- 0
x"00020",-- 2
x"000c0",-- 12
x"00080",-- 8
x"00000",-- 0
x"fffb0",-- -5
x"fffb0",-- -5
x"00000",-- 0
x"00030",-- 3
x"00000",-- 0
x"fffe0",-- -2
x"00000",-- 0
x"00000",-- 0
x"00020",-- 2
x"fffe0",-- -2
x"00000",-- 0
x"000d0",-- 13
x"00120",-- 18
x"00120",-- 18
x"00080",-- 8
x"000c0",-- 12
x"00080",-- 8
x"00080",-- 8
x"000a0",-- 10
x"00080",-- 8
x"00120",-- 18
x"00080",-- 8
x"00000",-- 0
x"00000",-- 0
x"fffb0",-- -5
x"00000",-- 0
x"fff60",-- -10
x"fff80",-- -8
x"00000",-- 0
x"fff10",-- -15
x"fff60",-- -10
x"00000",-- 0
x"fff40",-- -12
x"fffe0",-- -2
x"fffb0",-- -5
x"fff90",-- -7
x"fff60",-- -10
x"fffd0",-- -3
x"fffe0",-- -2
x"fffb0",-- -5
x"00000",-- 0
x"fff60",-- -10
x"fff30",-- -13
x"fff30",-- -13
x"fff90",-- -7
x"fff80",-- -8
x"fff90",-- -7
x"fff40",-- -12
x"ffef0",-- -17
x"ffea0",-- -22
x"fff10",-- -15
x"fff30",-- -13
x"ffec0",-- -20
x"fff10",-- -15
x"ffef0",-- -17
x"ffee0",-- -18
x"ffe40",-- -28
x"ffea0",-- -22
x"ffee0",-- -18
x"ffe70",-- -25
x"ffea0",-- -22
x"fff10",-- -15
x"ffdb0",-- -37
x"ffe50",-- -27
x"ffef0",-- -17
x"ffee0",-- -18
x"ffe70",-- -25
x"ffef0",-- -17
x"fff80",-- -8
x"ffe50",-- -27
x"ffe20",-- -30
x"ffe20",-- -30
x"ffdf0",-- -33
x"ffdb0",-- -37
x"ffd60",-- -42
x"ffd10",-- -47
x"ffc60",-- -58
x"ffda0",-- -38
x"ffd50",-- -43
x"ffd60",-- -42
x"ffdb0",-- -37
x"ffdf0",-- -33
x"ffd30",-- -45
x"ffc90",-- -55
x"ffc20",-- -62
x"ffc90",-- -55
x"ffb20",-- -78
x"fd850",-- -635
x"fbee0",-- -1042
x"fe0d0",-- -499
x"00c50",-- 197
x"ffa90",-- -87
x"ff010",-- -255
x"00e80",-- 232
x"021b0",-- 539
x"01ef0",-- 495
x"01770",-- 375
x"00530",-- 83
x"ff070",-- -249
x"ff600",-- -160
x"ff810",-- -127
x"ff8a0",-- -118
x"00460",-- 70
x"00ac0",-- 172
x"ffea0",-- -22
x"ffd10",-- -47
x"00a50",-- 165
x"fd900",-- -624
x"f9cc0",-- -1588
x"faf50",-- -1291
x"fe050",-- -507
x"fd4f0",-- -689
x"fd240",-- -732
x"ffd80",-- -40
x"017e0",-- 382
x"02dc0",-- 732
x"03330",-- 819
x"02260",-- 550
x"00850",-- 133
x"006c0",-- 108
x"ffb30",-- -77
x"ff350",-- -203
x"00460",-- 70
x"00760",-- 118
x"ffb50",-- -75
x"ff850",-- -123
x"00cd0",-- 205
x"ff810",-- -127
x"fe760",-- -394
x"fa660",-- -1434
x"ef720",-- -4238
x"eac80",-- -5432
x"f2a20",-- -3422
x"fce90",-- -791
x"01f40",-- 500
x"07450",-- 1861
x"0acf0",-- 2767
x"0ef00",-- 3824
x"10be0",-- 4286
x"0c810",-- 3201
x"02eb0",-- 747
x"fa170",-- -1513
x"f7400",-- -2240
x"f7d10",-- -2095
x"fc550",-- -939
x"015e0",-- 350
x"03ea0",-- 1002
x"03240",-- 804
x"040d0",-- 1037
x"03d10",-- 977
x"ffe40",-- -28
x"fa4d0",-- -1459
x"f5c00",-- -2624
x"f5a10",-- -2655
x"f8ed0",-- -1811
x"fe0a0",-- -502
x"00ff0",-- 255
x"03920",-- 914
x"06cd0",-- 1741
x"08b80",-- 2232
x"07770",-- 1911
x"051c0",-- 1308
x"02a00",-- 672
x"ffb00",-- -80
x"fe8c0",-- -372
x"ff130",-- -237
x"00110",-- 17
x"00190",-- 25
x"002f0",-- 47
x"001b0",-- 27
x"ff4a0",-- -182
x"fe980",-- -360
x"fcd00",-- -816
x"fa840",-- -1404
x"fa2b0",-- -1493
x"fbc10",-- -1087
x"fd710",-- -655
x"ffd80",-- -40
x"029d0",-- 669
x"046c0",-- 1132
x"055e0",-- 1374
x"05720",-- 1394
x"041b0",-- 1051
x"01810",-- 385
x"ffc60",-- -58
x"fe570",-- -425
x"fd200",-- -736
x"fd990",-- -615
x"ff1c0",-- -228
x"fff30",-- -13
x"00c80",-- 200
x"018f0",-- 399
x"00ed0",-- 237
x"00410",-- 65
x"ffdf0",-- -33
x"fef70",-- -265
x"fe660",-- -410
x"ff090",-- -247
x"ffee0",-- -18
x"00570",-- 87
x"01860",-- 390
x"025f0",-- 607
x"02520",-- 594
x"01ec0",-- 492
x"01810",-- 385
x"011f0",-- 287
x"010d0",-- 269
x"013f0",-- 319
x"01350",-- 309
x"01680",-- 360
x"02390",-- 569
x"025a0",-- 602
x"02190",-- 537
x"02490",-- 585
x"02260",-- 550
x"01380",-- 312
x"00df0",-- 223
x"01080",-- 264
x"01310",-- 305
x"00ac0",-- 172
x"009b0",-- 155
x"01090",-- 265
x"019a0",-- 410
x"02110",-- 529
x"01d00",-- 464
x"01d60",-- 470
x"01f60",-- 502
x"025c0",-- 604
x"020c0",-- 524
x"02800",-- 640
x"02750",-- 629
x"02990",-- 665
x"02aa0",-- 682
x"02b20",-- 690
x"02850",-- 645
x"01f10",-- 497
x"01650",-- 357
x"009b0",-- 155
x"00660",-- 102
x"00140",-- 20
x"ffad0",-- -83
x"ff790",-- -135
x"00300",-- 48
x"00a00",-- 160
x"00910",-- 145
x"00d90",-- 217
x"01450",-- 325
x"01180",-- 280
x"00230",-- 35
x"00080",-- 8
x"ff790",-- -135
x"fe170",-- -489
x"fcde0",-- -802
x"fc2d0",-- -979
x"fbc90",-- -1079
x"fb880",-- -1144
x"fbb00",-- -1104
x"fbbd0",-- -1091
x"fcbe0",-- -834
x"fd7e0",-- -642
x"fd7c0",-- -644
x"fd850",-- -635
x"fddf0",-- -545
x"fdf80",-- -520
x"fd1f0",-- -737
x"fce60",-- -794
x"fcad0",-- -851
x"fc390",-- -967
x"fbb70",-- -1097
x"fba90",-- -1111
x"fbf90",-- -1031
x"fc2b0",-- -981
x"fc6e0",-- -914
x"fc340",-- -972
x"fc8e0",-- -882
x"fd360",-- -714
x"fd5d0",-- -675
x"fd1b0",-- -741
x"fd490",-- -695
x"fd850",-- -635
x"fd4e0",-- -690
x"fd8a0",-- -630
x"fddb0",-- -549
x"fdc10",-- -575
x"fd760",-- -650
x"fe000",-- -512
x"fe7f0",-- -385
x"ff530",-- -173
x"fffb0",-- -5
x"ffea0",-- -22
x"00120",-- 18
x"00ac0",-- 172
x"01180",-- 280
x"00af0",-- 175
x"00490",-- 73
x"00200",-- 32
x"006c0",-- 108
x"00c80",-- 200
x"01740",-- 372
x"02120",-- 530
x"02890",-- 649
x"03fe0",-- 1022
x"05440",-- 1348
x"065d0",-- 1629
x"073d0",-- 1853
x"08580",-- 2136
x"091d0",-- 2333
x"08f20",-- 2290
x"08f90",-- 2297
x"08e60",-- 2278
x"08ff0",-- 2303
x"09650",-- 2405
x"0a930",-- 2707
x"0b0d0",-- 2829
x"0b880",-- 2952
x"0cca0",-- 3274
x"0d240",-- 3364
x"0d0b0",-- 3339
x"0bd00",-- 3024
x"0ae80",-- 2792
x"0ad20",-- 2770
x"0d120",-- 3346
x"0e930",-- 3731
x"0c7f0",-- 3199
x"088e0",-- 2190
x"040d0",-- 1037
x"fda10",-- -607
x"f47f0",-- -2945
x"ede00",-- -4640
x"e92f0",-- -5841
x"e6a50",-- -6491
x"e83a0",-- -6086
x"ee140",-- -4588
x"f5310",-- -2767
x"fc1e0",-- -994
x"00230",-- 35
x"016c0",-- 364
x"02e30",-- 739
x"02190",-- 537
x"ff150",-- -235
x"fbe50",-- -1051
x"fbba0",-- -1094
x"fc9e0",-- -866
x"fdea0",-- -534
x"ff720",-- -142
x"004d0",-- 77
x"ffa10",-- -95
x"fd3d0",-- -707
x"f9e20",-- -1566
x"f4eb0",-- -2837
x"f0e80",-- -3864
x"ed9a0",-- -4710
x"ec000",-- -5120
x"ed010",-- -4863
x"f0080",-- -4088
x"f3d60",-- -3114
x"f73e0",-- -2242
x"fabc0",-- -1348
x"fdbf0",-- -577
x"ff5b0",-- -165
x"ff440",-- -188
x"fea50",-- -347
x"fe2b0",-- -469
x"fe530",-- -429
x"fed40",-- -300
x"ff220",-- -222
x"ff380",-- -200
x"ff2b0",-- -213
x"fe930",-- -365
x"fd290",-- -727
x"fb070",-- -1273
x"f9200",-- -1760
x"f7ae0",-- -2130
x"f6e60",-- -2330
x"f79c0",-- -2148
x"f91d0",-- -1763
x"fb790",-- -1159
x"fe820",-- -382
x"01090",-- 265
x"03130",-- 787
x"049b0",-- 1179
x"05590",-- 1369
x"05150",-- 1301
x"04800",-- 1152
x"05060",-- 1286
x"05650",-- 1381
x"059c0",-- 1436
x"04c30",-- 1219
x"03cc0",-- 972
x"03620",-- 866
x"03d10",-- 977
x"03f40",-- 1012
x"03080",-- 776
x"02e60",-- 742
x"03210",-- 801
x"048e0",-- 1166
x"05950",-- 1429
x"06ac0",-- 1708
x"06b60",-- 1718
x"06f40",-- 1780
x"07ea0",-- 2026
x"097e0",-- 2430
x"0acc0",-- 2764
x"0af20",-- 2802
x"09f10",-- 2545
x"09d80",-- 2520
x"0be40",-- 3044
x"0ddf0",-- 3551
x"0f990",-- 3993
x"0f450",-- 3909
x"0ec80",-- 3784
x"10140",-- 4116
x"11bf0",-- 4543
x"0ff80",-- 4088
x"0cf20",-- 3314
x"0abe0",-- 2750
x"0aeb0",-- 2795
x"0ae30",-- 2787
x"091a0",-- 2330
x"04840",-- 1156
x"01bd0",-- 445
x"fff80",-- -8
x"fd830",-- -637
x"f7c70",-- -2105
x"f1900",-- -3696
x"eeac0",-- -4436
x"eeda0",-- -4390
x"f05c0",-- -4004
x"f1950",-- -3691
x"f6340",-- -2508
x"facf0",-- -1329
x"ff220",-- -222
x"01db0",-- 475
x"042f0",-- 1071
x"04b30",-- 1203
x"03810",-- 897
x"007f0",-- 127
x"feac0",-- -340
x"fe660",-- -410
x"fd1a0",-- -742
x"faca0",-- -1334
x"f9a40",-- -1628
x"fa8e0",-- -1394
x"f9970",-- -1641
x"f7ce0",-- -2098
x"f5ac0",-- -2644
x"f4c80",-- -2872
x"f3680",-- -3224
x"f2840",-- -3452
x"f2050",-- -3579
x"f2f00",-- -3344
x"f4ff0",-- -2817
x"f7040",-- -2300
x"f9450",-- -1723
x"fbba0",-- -1094
x"fe260",-- -474
x"feb20",-- -334
x"fec80",-- -312
x"ff4c0",-- -180
x"ffa30",-- -93
x"fec00",-- -320
x"fe370",-- -457
x"fd920",-- -622
x"fd3d0",-- -707
x"fcb70",-- -841
x"fbd80",-- -1064
x"fab10",-- -1359
x"f98b0",-- -1653
x"f8e30",-- -1821
x"f85d0",-- -1955
x"f8c10",-- -1855
x"f9b00",-- -1616
x"fb070",-- -1273
x"fcd50",-- -811
x"ffad0",-- -83
x"024b0",-- 587
x"03970",-- 919
x"04280",-- 1064
x"043c0",-- 1084
x"03f40",-- 1012
x"03600",-- 864
x"02390",-- 569
x"00750",-- 117
x"ff0b0",-- -245
x"ff7c0",-- -132
x"011f0",-- 287
x"02910",-- 657
x"039e0",-- 926
x"046e0",-- 1134
x"04ef0",-- 1263
x"05670",-- 1383
x"05ef0",-- 1519
x"056f0",-- 1391
x"04820",-- 1154
x"03c40",-- 964
x"04170",-- 1047
x"053a0",-- 1338
x"06ef0",-- 1775
x"086b0",-- 2155
x"09400",-- 2368
x"0afc0",-- 2812
x"0d150",-- 3349
x"0ec20",-- 3778
x"0fad0",-- 4013
x"10450",-- 4165
x"0f4c0",-- 3916
x"0dda0",-- 3546
x"0d1f0",-- 3359
x"0d220",-- 3362
x"0e0c0",-- 3596
x"0f330",-- 3891
x"0f680",-- 3944
x"0fb00",-- 4016
x"10f70",-- 4343
x"11090",-- 4361
x"0e640",-- 3684
x"0a780",-- 2680
x"07cb0",-- 1995
x"02210",-- 545
x"fa3f0",-- -1473
x"f3900",-- -3184
x"efdd0",-- -4131
x"eb790",-- -5255
x"e8690",-- -6039
x"ea350",-- -5579
x"eed00",-- -4400
x"f4670",-- -2969
x"f9160",-- -1770
x"fd850",-- -635
x"007a0",-- 122
x"02030",-- 515
x"008e0",-- 142
x"fe780",-- -392
x"fd440",-- -700
x"fc190",-- -999
x"fb0c0",-- -1268
x"fbb00",-- -1104
x"fd360",-- -714
x"fe210",-- -479
x"fdb20",-- -590
x"fbee0",-- -1042
x"fa390",-- -1479
x"f76d0",-- -2195
x"f4260",-- -3034
x"f0f00",-- -3856
x"ef650",-- -4251
x"eee60",-- -4378
x"ef6d0",-- -4243
x"f0760",-- -3978
x"f2930",-- -3437
x"f57e0",-- -2690
x"f7980",-- -2152
x"f94c0",-- -1716
x"faf20",-- -1294
x"fc7d0",-- -899
x"fd490",-- -695
x"fdf10",-- -527
x"fea80",-- -344
x"ff180",-- -232
x"ff130",-- -237
x"fed00",-- -304
x"fe230",-- -477
x"fce30",-- -797
x"fb790",-- -1159
x"f9c60",-- -1594
x"f8250",-- -2011
x"f7380",-- -2248
x"f7250",-- -2267
x"f7590",-- -2215
x"f8570",-- -1961
x"faa00",-- -1376
x"fd0c0",-- -756
x"ff1d0",-- -227
x"00b70",-- 183
x"01e50",-- 485
x"02cf0",-- 719
x"03bd0",-- 957
x"03fe0",-- 1022
x"03710",-- 881
x"031d0",-- 797
x"03210",-- 801
x"02e50",-- 741
x"03540",-- 852
x"03830",-- 899
x"03170",-- 791
x"028e0",-- 654
x"02a00",-- 672
x"02e30",-- 739
x"03260",-- 806
x"036a0",-- 874
x"03790",-- 889
x"04030",-- 1027
x"04850",-- 1157
x"056a0",-- 1386
x"05f10",-- 1521
x"07670",-- 1895
x"093a0",-- 2362
x"0b1d0",-- 2845
x"0d120",-- 3346
x"0ee60",-- 3814
x"0fcb0",-- 4043
x"10af0",-- 4271
x"10f40",-- 4340
x"0ff30",-- 4083
x"0df10",-- 3569
x"0bbf0",-- 3007
x"0b1a0",-- 2842
x"0b720",-- 2930
x"0d1c0",-- 3356
x"0f990",-- 3993
x"12c50",-- 4805
x"15360",-- 5430
x"15730",-- 5491
x"13f00",-- 5104
x"11470",-- 4423
x"0d2e0",-- 3374
x"083f0",-- 2111
x"030d0",-- 781
x"fe210",-- -479
x"f8390",-- -1991
x"f2f80",-- -3336
x"ef480",-- -4280
x"ee210",-- -4575
x"ee700",-- -4496
x"ee2e0",-- -4562
x"eeb10",-- -4431
x"f1fb0",-- -3589
x"f6d90",-- -2343
x"f90b0",-- -1781
x"fa210",-- -1503
x"fb5b0",-- -1189
x"fc3f0",-- -961
x"fd1b0",-- -741
x"fe1c0",-- -484
x"fefd0",-- -259
x"00840",-- 132
x"01a10",-- 417
x"01c20",-- 450
x"01ce0",-- 462
x"00c50",-- 197
x"fdfd0",-- -515
x"f9e90",-- -1559
x"f67b0",-- -2437
x"f2e40",-- -3356
x"efab0",-- -4181
x"ed1b0",-- -4837
x"ebb10",-- -5199
x"ebb30",-- -5197
x"ece30",-- -4893
x"eed40",-- -4396
x"f11a0",-- -3814
x"f51d0",-- -2787
x"f8c80",-- -1848
x"fbb70",-- -1097
x"fea50",-- -347
x"01130",-- 275
x"02760",-- 630
x"02d40",-- 724
x"02350",-- 565
x"00af0",-- 175
x"fea50",-- -347
x"fc870",-- -889
x"fa990",-- -1383
x"f8f70",-- -1801
x"f7ae0",-- -2130
x"f6690",-- -2455
x"f62f0",-- -2513
x"f72f0",-- -2257
x"f83f0",-- -1985
x"f9a90",-- -1623
x"fb6c0",-- -1172
x"fd5d0",-- -675
x"fef80",-- -264
x"007a0",-- 122
x"018a0",-- 394
x"02620",-- 610
x"03330",-- 819
x"03810",-- 897
x"03cc0",-- 972
x"03c70",-- 967
x"04480",-- 1096
x"04be0",-- 1214
x"05240",-- 1316
x"05920",-- 1426
x"05720",-- 1394
x"056f0",-- 1391
x"055e0",-- 1374
x"04f00",-- 1264
x"03ec0",-- 1004
x"02ed0",-- 749
x"01c20",-- 450
x"014e0",-- 334
x"019e0",-- 414
x"02f40",-- 756
x"04800",-- 1152
x"066c0",-- 1644
x"08ea0",-- 2282
x"0b580",-- 2904
x"0da80",-- 3496
x"0eb40",-- 3764
x"0f350",-- 3893
x"0f010",-- 3841
x"0e930",-- 3731
x"0dbd0",-- 3517
x"0d2e0",-- 3374
x"0cca0",-- 3274
x"0b800",-- 2944
x"0ab30",-- 2739
x"0b7c0",-- 2940
x"0df50",-- 3573
x"0f800",-- 3968
x"10950",-- 4245
x"12540",-- 4692
x"14310",-- 5169
x"13b00",-- 5040
x"117e0",-- 4478
x"0f1f0",-- 3871
x"0d4c0",-- 3404
x"09950",-- 2453
x"03530",-- 851
x"fc3f0",-- -961
x"f72e0",-- -2258
x"f5a70",-- -2649
x"f1d30",-- -3629
x"ece60",-- -4890
x"ea8a0",-- -5494
x"ec820",-- -4990
x"ee870",-- -4473
x"f08c0",-- -3956
x"f2640",-- -3484
x"f4480",-- -3000
x"f6490",-- -2487
x"f7950",-- -2155
x"fa710",-- -1423
x"fd330",-- -717
x"ff270",-- -217
x"ff920",-- -110
x"01150",-- 277
x"03b00",-- 944
x"04c00",-- 1216
x"02ed0",-- 749
x"ff760",-- -138
x"fc1c0",-- -996
x"f9070",-- -1785
x"f5180",-- -2792
x"f02b0",-- -4053
x"eca20",-- -4958
x"ead20",-- -5422
x"e9d80",-- -5672
x"ea2d0",-- -5587
x"ec440",-- -5052
x"eef70",-- -4361
x"f1e00",-- -3616
x"f5160",-- -2794
x"f9070",-- -1785
x"fcaa0",-- -854
x"fec80",-- -312
x"00110",-- 17
x"00e40",-- 228
x"014f0",-- 335
x"01180",-- 280
x"003a0",-- 58
x"fefa0",-- -262
x"fd8a0",-- -630
x"fc260",-- -986
x"fad40",-- -1324
x"f9c10",-- -1599
x"f8b70",-- -1865
x"f7b50",-- -2123
x"f7520",-- -2222
x"f7ba0",-- -2118
x"f8da0",-- -1830
x"fa320",-- -1486
x"fb240",-- -1244
x"fca20",-- -862
x"fe910",-- -367
x"008c0",-- 140
x"02250",-- 549
x"039e0",-- 926
x"04c50",-- 1221
x"053d0",-- 1341
x"05e40",-- 1508
x"061b0",-- 1563
x"06300",-- 1584
x"05ce0",-- 1486
x"05830",-- 1411
x"05720",-- 1394
x"05a80",-- 1448
x"061e0",-- 1566
x"06110",-- 1553
x"05860",-- 1414
x"053b0",-- 1339
x"04990",-- 1177
x"03740",-- 884
x"029e0",-- 670
x"02db0",-- 731
x"03fe0",-- 1022
x"051d0",-- 1309
x"06ff0",-- 1791
x"08ff0",-- 2303
x"0ae80",-- 2792
x"0c020",-- 3074
x"0c810",-- 3201
x"0ccf0",-- 3279
x"0ccc0",-- 3276
x"0cd20",-- 3282
x"0cc50",-- 3269
x"0ca50",-- 3237
x"0cdc0",-- 3292
x"0cf50",-- 3317
x"0dda0",-- 3546
x"0e5a0",-- 3674
x"0f3a0",-- 3898
x"10ef0",-- 4335
x"130d0",-- 4877
x"14250",-- 5157
x"13bf0",-- 5055
x"13180",-- 4888
x"123e0",-- 4670
x"10630",-- 4195
x"0d800",-- 3456
x"0bd60",-- 3030
x"08ef0",-- 2287
x"031c0",-- 796
x"fc390",-- -967
x"f84e0",-- -1970
x"f4750",-- -2955
x"ee850",-- -4475
x"e88a0",-- -6006
x"e6d80",-- -6440
x"e8050",-- -6139
x"e9740",-- -5772
x"ec4c0",-- -5044
x"f12a0",-- -3798
x"f6250",-- -2523
x"f9340",-- -1740
x"fc370",-- -969
x"ff1f0",-- -225
x"01a40",-- 420
x"022b0",-- 555
x"01540",-- 340
x"00b20",-- 178
x"01a40",-- 420
x"01580",-- 344
x"ff010",-- -255
x"fcaa0",-- -854
x"fae90",-- -1303
x"f7d80",-- -2088
x"f4210",-- -3039
x"f1950",-- -3691
x"efab0",-- -4181
x"ed470",-- -4793
x"eb150",-- -5355
x"eb4c0",-- -5300
x"ed360",-- -4810
x"ef6a0",-- -4246
x"f15e0",-- -3746
x"f45d0",-- -2979
x"f80d0",-- -2035
x"fba10",-- -1119
x"fe120",-- -494
x"ffd00",-- -48
x"00eb0",-- 235
x"01380",-- 312
x"007d0",-- 125
x"ffee0",-- -18
x"ffa60",-- -90
x"febb0",-- -325
x"fcff0",-- -769
x"fb9a0",-- -1126
x"fb5e0",-- -1186
x"fafd0",-- -1283
x"fa030",-- -1533
x"f8fc0",-- -1796
x"f8ad0",-- -1875
x"f8b70",-- -1865
x"f9380",-- -1736
x"fa390",-- -1479
x"fbf80",-- -1032
x"fdc10",-- -575
x"ff630",-- -157
x"01580",-- 344
x"03ba0",-- 954
x"05600",-- 1376
x"05ce0",-- 1486
x"05ec0",-- 1516
x"067a0",-- 1658
x"07090",-- 1801
x"071d0",-- 1821
x"07440",-- 1860
x"07880",-- 1928
x"07fb0",-- 2043
x"07ea0",-- 2026
x"07770",-- 1911
x"06d90",-- 1753
x"05cc0",-- 1484
x"04610",-- 1121
x"03040",-- 772
x"02730",-- 627
x"02250",-- 549
x"023c0",-- 572
x"02bc0",-- 700
x"04000",-- 1024
x"060f0",-- 1551
x"07dd0",-- 2013
x"097e0",-- 2430
x"0aaa0",-- 2730
x"0bbf0",-- 3007
x"0c6d0",-- 3181
x"0cd70",-- 3287
x"0d2b0",-- 3371
x"0d4c0",-- 3404
x"0d270",-- 3367
x"0d470",-- 3399
x"0dbc0",-- 3516
x"0e230",-- 3619
x"0ec30",-- 3779
x"104b0",-- 4171
x"12b60",-- 4790
x"14090",-- 5129
x"147c0",-- 5244
x"14930",-- 5267
x"13f50",-- 5109
x"12310",-- 4657
x"0f0d0",-- 3853
x"0c7c0",-- 3196
x"091a0",-- 2330
x"037b0",-- 891
x"fc780",-- -904
x"f71d0",-- -2275
x"f32a0",-- -3286
x"ee7d0",-- -4483
x"ea8a0",-- -5494
x"e7790",-- -6279
x"e7bd0",-- -6211
x"e9fc0",-- -5636
x"ec5b0",-- -5029
x"eeed0",-- -4371
x"f28c0",-- -3444
x"f58e0",-- -2674
x"f7930",-- -2157
x"f9dd0",-- -1571
x"fc760",-- -906
x"fe890",-- -375
x"ff130",-- -237
x"fffb0",-- -5
x"01a90",-- 425
x"03740",-- 884
x"037b0",-- 891
x"03210",-- 801
x"01ce0",-- 462
x"ff970",-- -105
x"fc4e0",-- -946
x"f7950",-- -2155
x"f3270",-- -3289
x"efea0",-- -4118
x"ecbc0",-- -4932
x"e9610",-- -5791
x"e8d20",-- -5934
x"ea290",-- -5591
x"ec6a0",-- -5014
x"eefc0",-- -4356
x"f2d20",-- -3374
x"f7130",-- -2285
x"fa990",-- -1383
x"fd270",-- -729
x"ff6d0",-- -147
x"013f0",-- 319
x"01cc0",-- 460
x"01b30",-- 435
x"011a0",-- 282
x"00cf0",-- 207
x"00760",-- 118
x"ffad0",-- -83
x"fee30",-- -285
x"fead0",-- -339
x"fde00",-- -544
x"fc990",-- -871
x"fb710",-- -1167
x"fac10",-- -1343
x"fa2b0",-- -1493
x"f97c0",-- -1668
x"f9bf0",-- -1601
x"faad0",-- -1363
x"fc1c0",-- -996
x"fe030",-- -509
x"00800",-- 128
x"03330",-- 819
x"05600",-- 1376
x"06d10",-- 1745
x"07a30",-- 1955
x"088e0",-- 2190
x"09310",-- 2353
x"08f40",-- 2292
x"080f0",-- 2063
x"077b0",-- 1915
x"06f50",-- 1781
x"06320",-- 1586
x"05b70",-- 1463
x"05510",-- 1361
x"04800",-- 1152
x"03240",-- 804
x"02480",-- 584
x"01c20",-- 450
x"01540",-- 340
x"00fc0",-- 252
x"00ff0",-- 255
x"01ce0",-- 462
x"034a0",-- 842
x"05150",-- 1301
x"06d10",-- 1745
x"08840",-- 2180
x"0a450",-- 2629
x"0b650",-- 2917
x"0bf40",-- 3060
x"0c3e0",-- 3134
x"0c3e0",-- 3134
x"0bb30",-- 2995
x"0b0d0",-- 2829
x"0acc0",-- 2764
x"0afe0",-- 2814
x"0b530",-- 2899
x"0bbc0",-- 3004
x"0c3b0",-- 3131
x"0cc80",-- 3272
x"0dae0",-- 3502
x"0ea50",-- 3749
x"0f990",-- 3993
x"0fa10",-- 4001
x"0f0e0",-- 3854
x"0de70",-- 3559
x"0d7b0",-- 3451
x"0c0d0",-- 3085
x"09130",-- 2323
x"05080",-- 1288
x"01060",-- 262
x"fce80",-- -792
x"f8410",-- -1983
x"f4550",-- -2987
x"f0a20",-- -3934
x"edfc0",-- -4612
x"ec030",-- -5117
x"ebcc0",-- -5172
x"ecb90",-- -4935
x"ee7a0",-- -4486
x"f0190",-- -4071
x"f1920",-- -3694
x"f3660",-- -3226
x"f59a0",-- -2662
x"f7740",-- -2188
x"f8a20",-- -1886
x"f9f80",-- -1544
x"fb5e0",-- -1186
x"fcf00",-- -784
x"fe210",-- -479
x"ffe20",-- -30
x"01420",-- 322
x"019e0",-- 414
x"00d00",-- 208
x"00000",-- 0
x"fedf0",-- -289
x"fcfd0",-- -771
x"fa350",-- -1483
x"f72c0",-- -2260
x"f5110",-- -2799
x"f39d0",-- -3171
x"f2bb0",-- -3397
x"f2620",-- -3486
x"f31f0",-- -3297
x"f4460",-- -3002
x"f58e0",-- -2674
x"f7430",-- -2237
x"f96d0",-- -1683
x"fb360",-- -1226
x"fbf90",-- -1031
x"fc260",-- -986
x"fc820",-- -894
x"fcf00",-- -784
x"fd110",-- -751
x"fced0",-- -787
x"fcb20",-- -846
x"fcc60",-- -826
x"fd270",-- -729
x"fd920",-- -622
x"fe370",-- -457
x"ff2e0",-- -210
x"ffc40",-- -60
x"00250",-- 37
x"00f00",-- 240
x"02210",-- 545
x"033a0",-- 826
x"03cc0",-- 972
x"04490",-- 1097
x"04e10",-- 1249
x"05770",-- 1399
x"05da0",-- 1498
x"05fb0",-- 1531
x"05e90",-- 1513
x"05a30",-- 1443
x"052c0",-- 1324
x"04990",-- 1177
x"04140",-- 1044
x"03a10",-- 929
x"03080",-- 776
x"02750",-- 629
x"01fe0",-- 510
x"01dd0",-- 477
x"019a0",-- 410
x"01420",-- 322
x"01180",-- 280
x"00ef0",-- 239
x"00ef0",-- 239
x"00cf0",-- 207
x"00e80",-- 232
x"014e0",-- 334
x"01b30",-- 435
x"02320",-- 562
x"02e10",-- 737
x"03490",-- 841
x"039e0",-- 926
x"03f40",-- 1012
x"03ee0",-- 1006
x"03d10",-- 977
x"03c90",-- 969
x"037c0",-- 892
x"03100",-- 784
x"02ca0",-- 714
x"02640",-- 612
x"021b0",-- 539
x"01d00",-- 464
x"01a40",-- 420
x"01db0",-- 475
x"02030",-- 515
x"025c0",-- 604
x"02fe0",-- 766
x"039a0",-- 922
x"042a0",-- 1066
x"04b30",-- 1203
x"05490",-- 1353
x"061e0",-- 1566
x"06c80",-- 1736
x"073b0",-- 1851
x"078f0",-- 1935
x"07dd0",-- 2013
x"080c0",-- 2060
x"07d30",-- 2003
x"07470",-- 1863
x"06960",-- 1686
x"06070",-- 1543
x"054a0",-- 1354
x"042d0",-- 1069
x"03380",-- 824
x"02610",-- 609
x"01620",-- 354
x"00430",-- 67
x"ff600",-- -160
x"fea00",-- -352
x"fd990",-- -615
x"fc7a0",-- -902
x"fb650",-- -1179
x"fa480",-- -1464
x"f92f0",-- -1745
x"f8390",-- -1991
x"f73e0",-- -2242
x"f6af0",-- -2385
x"f6a20",-- -2398
x"f6e80",-- -2328
x"f78e0",-- -2162
x"f8a50",-- -1883
x"f9df0",-- -1569
x"fae80",-- -1304
x"fbbd0",-- -1091
x"fc6b0",-- -917
x"fced0",-- -787
x"fd020",-- -766
x"fcd50",-- -811
x"fc8f0",-- -881
x"fc260",-- -986
x"fbd00",-- -1072
x"fb8b0",-- -1141
x"fb420",-- -1214
x"fafa0",-- -1286
x"fac60",-- -1338
x"fac60",-- -1338
x"fad90",-- -1319
x"fadf0",-- -1313
x"facf0",-- -1329
x"fac80",-- -1336
x"fa8a0",-- -1398
x"fa6e0",-- -1426
x"fa3e0",-- -1474
x"fa3e0",-- -1474
x"fa7f0",-- -1409
x"fadf0",-- -1313
x"fb5c0",-- -1188
x"fc190",-- -999
x"fd2c0",-- -724
x"fe640",-- -412
x"ff970",-- -105
x"00b40",-- 180
x"01b70",-- 439
x"02890",-- 649
x"03650",-- 869
x"03e50",-- 997
x"04250",-- 1061
x"043f0",-- 1087
x"04460",-- 1094
x"04230",-- 1059
x"03e40",-- 996
x"03a80",-- 936
x"03760",-- 886
x"03450",-- 837
x"02eb0",-- 747
x"02b20",-- 690
x"027a0",-- 634
x"02260",-- 550
x"01db0",-- 475
x"018a0",-- 394
x"01360",-- 310
x"01120",-- 274
x"01120",-- 274
x"01180",-- 280
x"01210",-- 289
x"014f0",-- 335
x"01c20",-- 450
x"01fd0",-- 509
x"02230",-- 547
x"02500",-- 592
x"02500",-- 592
x"022b0",-- 555
x"01e40",-- 484
x"018d0",-- 397
x"01180",-- 280
x"00b60",-- 182
x"00570",-- 87
x"00000",-- 0
x"ffbf0",-- -65
x"ffa90",-- -87
x"ff900",-- -112
x"ff920",-- -110
x"ffab0",-- -85
x"ffa30",-- -93
x"ffb50",-- -75
x"ffb30",-- -77
x"ff9f0",-- -97
x"ff830",-- -125
x"ff6d0",-- -147
x"ff330",-- -205
x"ff270",-- -217
x"ff110",-- -239
x"ff260",-- -218
x"ff6a0",-- -150
x"ffbd0",-- -67
x"00430",-- 67
x"00c50",-- 197
x"01530",-- 339
x"01d30",-- 467
x"02640",-- 612
x"02ea0",-- 746
x"03680",-- 872
x"03e50",-- 997
x"04640",-- 1124
x"04f00",-- 1264
x"055e0",-- 1374
x"05ba0",-- 1466
x"05bd0",-- 1469
x"058f0",-- 1423
x"055b0",-- 1371
x"05210",-- 1313
x"04c50",-- 1221
x"04350",-- 1077
x"03cb0",-- 971
x"03490",-- 841
x"02d40",-- 724
x"02980",-- 664
x"02690",-- 617
x"021e0",-- 542
x"01ce0",-- 462
x"01450",-- 325
x"00bc0",-- 188
x"00410",-- 65
x"ffb80",-- -72
x"ff100",-- -240
x"fe500",-- -432
x"fdb20",-- -590
x"fd340",-- -716
x"fce30",-- -797
x"fcaa0",-- -854
x"fc980",-- -872
x"fc910",-- -879
x"fc890",-- -887
x"fc8f0",-- -881
x"fca30",-- -861
x"fcb10",-- -847
x"fc9e0",-- -866
x"fc7f0",-- -897
x"fc3e0",-- -962
x"fc030",-- -1021
x"fbd50",-- -1067
x"fb940",-- -1132
x"fb590",-- -1191
x"fb1d0",-- -1251
x"faf50",-- -1291
x"fadc0",-- -1316
x"fb020",-- -1278
x"fb570",-- -1193
x"fb8d0",-- -1139
x"fbec0",-- -1044
x"fc620",-- -926
x"fcdc0",-- -804
x"fd580",-- -680
x"fdda0",-- -550
x"fe530",-- -429
x"fe9e0",-- -354
x"fed50",-- -299
x"fee90",-- -279
x"fee30",-- -285
x"fedf0",-- -289
x"fec30",-- -317
x"fea80",-- -344
x"fea70",-- -345
x"fee30",-- -285
x"ff300",-- -208
x"ff8a0",-- -118
x"fffb0",-- -5
x"005d0",-- 93
x"00cf0",-- 207
x"013b0",-- 315
x"01ba0",-- 442
x"022d0",-- 557
x"028e0",-- 654
x"02e10",-- 737
x"03180",-- 792
x"03330",-- 819
x"031f0",-- 799
x"02f50",-- 757
x"02ca0",-- 714
x"029d0",-- 669
x"02500",-- 592
x"020a0",-- 522
x"01e50",-- 485
x"01d00",-- 464
x"01d30",-- 467
x"01c10",-- 449
x"01b70",-- 439
x"01b70",-- 439
x"01ba0",-- 442
x"01b00",-- 432
x"01990",-- 409
x"016f0",-- 367
x"011d0",-- 285
x"00e30",-- 227
x"007d0",-- 125
x"001e0",-- 30
x"ffc20",-- -62
x"ff800",-- -128
x"ff440",-- -188
x"fefa0",-- -262
x"fef00",-- -272
x"fee30",-- -285
x"fee30",-- -285
x"fee60",-- -282
x"fef70",-- -265
x"ff220",-- -222
x"ff4a0",-- -182
x"ff830",-- -125
x"ffa30",-- -93
x"ffa90",-- -87
x"ffea0",-- -22
x"fff40",-- -12
x"ffd80",-- -40
x"fff10",-- -15
x"000c0",-- 12
x"001c0",-- 28
x"002a0",-- 42
x"006e0",-- 110
x"00b90",-- 185
x"00ef0",-- 239
x"01300",-- 304
x"01720",-- 370
x"01a60",-- 422
x"02020",-- 514
x"024b0",-- 587
x"02930",-- 659
x"03010",-- 769
x"036f0",-- 879
x"03d60",-- 982
x"04170",-- 1047
x"04780",-- 1144
x"04850",-- 1157
x"045f0",-- 1119
x"04410",-- 1089
x"04300",-- 1072
x"04050",-- 1029
x"03b00",-- 944
x"037b0",-- 891
x"03380",-- 824
x"02fe0",-- 766
x"02b40",-- 692
x"025f0",-- 607
x"02080",-- 520
x"01a10",-- 417
x"010e0",-- 270
x"00640",-- 100
x"ffe50",-- -27
x"ff540",-- -172
x"febb0",-- -325
x"fe200",-- -480
x"fda40",-- -604
x"fd510",-- -687
x"fd090",-- -759
x"fcdf0",-- -801
x"fcda0",-- -806
x"fcde0",-- -802
x"fce60",-- -794
x"fcdc0",-- -804
x"fcd40",-- -812
x"fcda0",-- -806
x"fcd50",-- -811
x"fc910",-- -879
x"fc4b0",-- -949
x"fc350",-- -971
x"fc050",-- -1019
x"fbdf0",-- -1057
x"fbc90",-- -1079
x"fbbf0",-- -1089
x"fbda0",-- -1062
x"fbdd0",-- -1059
x"fbf40",-- -1036
x"fc2d0",-- -979
x"fc550",-- -939
x"fc8f0",-- -881
x"fca70",-- -857
x"fcd70",-- -809
x"fd160",-- -746
x"fd360",-- -714
x"fd5d0",-- -675
x"fd6c0",-- -660
x"fd920",-- -622
x"fdb80",-- -584
x"fde40",-- -540
x"fe370",-- -457
x"fe820",-- -382
x"fec10",-- -319
x"ff170",-- -233
x"ff850",-- -123
x"fff80",-- -8
x"00690",-- 105
x"00d70",-- 215
x"013b0",-- 315
x"01a30",-- 419
x"01e50",-- 485
x"020a0",-- 522
x"02340",-- 564
x"02370",-- 567
x"02140",-- 532
x"01ef0",-- 495
x"01e20",-- 482
x"01df0",-- 479
x"01ce0",-- 462
x"01ba0",-- 442
x"019a0",-- 410
x"01a30",-- 419
x"01a30",-- 419
x"01b00",-- 432
x"01c10",-- 449
x"01d80",-- 472
x"01f10",-- 497
x"01c60",-- 454
x"01da0",-- 474
x"01a90",-- 425
x"018b0",-- 395
x"01830",-- 387
x"01490",-- 329
x"01180",-- 280
x"00eb0",-- 235
x"00be0",-- 190
x"00870",-- 135
x"00730",-- 115
x"00580",-- 88
x"00430",-- 67
x"00250",-- 37
x"000a0",-- 10
x"00120",-- 18
x"001e0",-- 30
x"00160",-- 22
x"00200",-- 32
x"00280",-- 40
x"00140",-- 20
x"002a0",-- 42
x"00370",-- 55
x"00370",-- 55
x"005a0",-- 90
x"008c0",-- 140
x"00af0",-- 175
x"00df0",-- 223
x"01240",-- 292
x"01790",-- 377
x"01c40",-- 452
x"020a0",-- 522
x"025d0",-- 605
x"028c0",-- 652
x"02bb0",-- 699
x"02ed0",-- 749
x"030d0",-- 781
x"03310",-- 817
x"032c0",-- 812
x"02f40",-- 756
x"02c60",-- 710
x"02ad0",-- 685
x"02750",-- 629
x"023f0",-- 575
x"02070",-- 519
x"01c60",-- 454
x"01a80",-- 424
x"017e0",-- 382
x"01540",-- 340
x"011f0",-- 287
x"00e40",-- 228
x"00800",-- 128
x"00140",-- 20
x"ffc90",-- -55
x"ff6c0",-- -148
x"fef30",-- -269
x"fe760",-- -394
x"fe030",-- -509
x"fd9c0",-- -612
x"fd4c0",-- -692
x"fd0c0",-- -756
x"fce90",-- -791
x"fcca0",-- -822
x"fcb40",-- -844
x"fc9e0",-- -866
x"fc8a0",-- -886
x"fc910",-- -879
x"fc940",-- -876
x"fc750",-- -907
x"fc5d0",-- -931
x"fc670",-- -921
x"fc5c0",-- -932
x"fc530",-- -941
x"fc460",-- -954
x"fc3c0",-- -964
x"fc3f0",-- -961
x"fc210",-- -991
x"fc170",-- -1001
x"fc320",-- -974
x"fc390",-- -967
x"fc460",-- -954
x"fc610",-- -927
x"fc6c0",-- -916
x"fcaa0",-- -854
x"fceb0",-- -789
x"fd330",-- -717
x"fd710",-- -655
x"fdb00",-- -592
x"fe080",-- -504
x"fe490",-- -439
x"fe9d0",-- -355
x"fede0",-- -290
x"ff150",-- -235
x"ff5d0",-- -163
x"ff850",-- -123
x"ffc40",-- -60
x"00170",-- 23
x"00520",-- 82
x"00990",-- 153
x"00d90",-- 217
x"010d0",-- 269
x"014a0",-- 330
x"01970",-- 407
x"01c90",-- 457
x"01e50",-- 485
x"01f90",-- 505
x"020d0",-- 525
x"02230",-- 547
x"022f0",-- 559
x"02490",-- 585
x"02440",-- 580
x"023c0",-- 572
x"02390",-- 569
x"021c0",-- 540
x"02080",-- 520
x"01fd0",-- 509
x"01fd0",-- 509
x"02020",-- 514
x"01e50",-- 485
x"01e70",-- 487
x"01d50",-- 469
x"01ba0",-- 442
x"01a30",-- 419
x"01830",-- 387
x"01620",-- 354
x"01270",-- 295
x"01080",-- 264
x"00c50",-- 197
x"009d0",-- 157
x"007d0",-- 125
x"00410",-- 65
x"003a0",-- 58
x"003c0",-- 60
x"00480",-- 72
x"004b0",-- 75
x"00480",-- 72
x"006e0",-- 110
x"00870",-- 135
x"00870",-- 135
x"008f0",-- 143
x"00a80",-- 168
x"00b20",-- 178
x"00b10",-- 177
x"00bc0",-- 188
x"00d20",-- 210
x"00ed0",-- 237
x"00f50",-- 245
x"01090",-- 265
x"01360",-- 310
x"01510",-- 337
x"01810",-- 385
x"01b50",-- 437
x"01f30",-- 499
x"022a0",-- 554
x"02690",-- 617
x"02a00",-- 672
x"02c00",-- 704
x"02bc0",-- 700
x"02ac0",-- 684
x"028f0",-- 655
x"026e0",-- 622
x"02410",-- 577
x"01f60",-- 502
x"01bf0",-- 447
x"018a0",-- 394
x"01560",-- 342
x"011f0",-- 287
x"00f50",-- 245
x"00c50",-- 197
x"00760",-- 118
x"00230",-- 35
x"ffc90",-- -55
x"ff7c0",-- -132
x"ff240",-- -220
x"fec60",-- -314
x"fe660",-- -410
x"fe170",-- -489
x"fdc60",-- -570
x"fd7c0",-- -644
x"fd470",-- -697
x"fd0e0",-- -754
x"fcfc0",-- -772
x"fced0",-- -787
x"fcc10",-- -831
x"fcb40",-- -844
x"fccd0",-- -819
x"fcb60",-- -842
x"fca50",-- -859
x"fc930",-- -877
x"fc980",-- -872
x"fca80",-- -856
x"fca50",-- -859
x"fcb70",-- -841
x"fcad0",-- -851
x"fc890",-- -887
x"fc9e0",-- -866
x"fcc30",-- -829
x"fcc60",-- -826
x"fcca0",-- -822
x"fcd70",-- -809
x"fcf80",-- -776
x"fd240",-- -732
x"fd2c0",-- -724
x"fd4f0",-- -689
x"fda10",-- -607
x"fdc10",-- -575
x"fdef0",-- -529
x"fe2d0",-- -467
x"fe870",-- -377
x"fec00",-- -320
x"ff0b0",-- -245
x"ff510",-- -175
x"ff8d0",-- -115
x"ffee0",-- -18
x"00160",-- 22
x"00760",-- 118
x"00990",-- 153
x"00d00",-- 208
x"00fa0",-- 250
x"01220",-- 290
x"01590",-- 345
x"01790",-- 377
x"019f0",-- 415
x"01a90",-- 425
x"01d30",-- 467
x"01e20",-- 482
x"01f30",-- 499
x"02000",-- 512
x"02070",-- 519
x"02070",-- 519
x"02020",-- 514
x"02000",-- 512
x"01f30",-- 499
x"01ef0",-- 495
x"01e40",-- 484
x"01d10",-- 465
x"01b50",-- 437
x"01ad0",-- 429
x"01b30",-- 435
x"01860",-- 390
x"016f0",-- 367
x"01590",-- 345
x"01450",-- 325
x"013f0",-- 319
x"01350",-- 309
x"01130",-- 275
x"00ed0",-- 237
x"00cf0",-- 207
x"00c00",-- 192
x"00ac0",-- 172
x"00800",-- 128
x"00730",-- 115
x"00660",-- 102
x"00710",-- 113
x"006b0",-- 107
x"00800",-- 128
x"00870",-- 135
x"00a30",-- 163
x"00bb0",-- 187
x"00d50",-- 213
x"00f70",-- 247
x"01090",-- 265
x"01260",-- 294
x"01310",-- 305
x"01560",-- 342
x"01620",-- 354
x"016f0",-- 367
x"019e0",-- 414
x"01b00",-- 432
x"01df0",-- 479
x"02250",-- 549
x"02460",-- 582
x"02660",-- 614
x"02910",-- 657
x"029d0",-- 669
x"02aa0",-- 682
x"02940",-- 660
x"027f0",-- 639
x"026b0",-- 619
x"02300",-- 560
x"01f90",-- 505
x"01bd0",-- 445
x"018a0",-- 394
x"013b0",-- 315
x"00f40",-- 244
x"00bb0",-- 187
x"00800",-- 128
x"002a0",-- 42
x"fff10",-- -15
x"ffa80",-- -88
x"ff170",-- -233
x"fefa0",-- -262
x"fe7f0",-- -385
x"fe300",-- -464
x"fe110",-- -495
x"fdab0",-- -597
x"fd7b0",-- -645
x"fd5b0",-- -677
x"fd400",-- -704
x"fd160",-- -746
x"fd530",-- -685
x"fd200",-- -736
x"fd0b0",-- -757
x"fd180",-- -744
x"fcf20",-- -782
x"fcd00",-- -816
x"fce90",-- -791
x"fcf70",-- -777
x"fcc60",-- -826
x"fcfc0",-- -772
x"fcd40",-- -812
x"fcda0",-- -806
x"fd1d0",-- -739
x"fd020",-- -766
x"fd2c0",-- -724
x"fd180",-- -744
x"fd160",-- -746
x"fd4c0",-- -692
x"fd560",-- -682
x"fd6f0",-- -657
x"fd850",-- -635
x"fd990",-- -615
x"fdab0",-- -597
x"fde50",-- -539
x"fe210",-- -479
x"fe6c0",-- -404
x"fee80",-- -280
x"ff010",-- -255
x"ff170",-- -233
x"ff5e0",-- -162
x"ffa10",-- -95
x"00020",-- 2
x"00660",-- 102
x"00c00",-- 192
x"00c50",-- 197
x"013d0",-- 317
x"015e0",-- 350
x"01380",-- 312
x"016a0",-- 362
x"017b0",-- 379
x"01cc0",-- 460
x"01a90",-- 425
x"01b70",-- 439
x"02050",-- 517
x"02340",-- 564
x"02480",-- 584
x"02520",-- 594
x"022f0",-- 559
x"02030",-- 515
x"017c0",-- 380
x"01ec0",-- 492
x"02000",-- 512
x"01fb0",-- 507
x"01bd0",-- 445
x"01b00",-- 432
x"01e90",-- 489
x"019e0",-- 414
x"01ce0",-- 462
x"016a0",-- 362
x"01470",-- 327
x"01800",-- 384
x"01060",-- 262
x"00a80",-- 168
x"01310",-- 305
x"016a0",-- 362
x"01680",-- 360
x"01450",-- 325
x"01760",-- 374
x"01970",-- 407
x"00f90",-- 249
x"00d20",-- 210
x"01260",-- 294
x"00cf0",-- 207
x"00d00",-- 208
x"00990",-- 153
x"00e80",-- 232
x"014e0",-- 334
x"01d10",-- 465
x"01400",-- 320
x"01e50",-- 485
x"02050",-- 517
x"01040",-- 260
x"02210",-- 545
x"014e0",-- 334
x"01f90",-- 505
x"02520",-- 594
x"02160",-- 534
x"029b0",-- 667
x"02a00",-- 672
x"034f0",-- 847
x"02d40",-- 724
x"02fe0",-- 766
x"02c80",-- 712
x"025c0",-- 604
x"02a70",-- 679
x"02520",-- 594
x"01e50",-- 485
x"01f30",-- 499
x"01860",-- 390
x"01720",-- 370
x"01560",-- 342
x"00910",-- 145
x"00990",-- 153
x"007f0",-- 127
x"ffbf0",-- -65
x"ff600",-- -160
x"ff540",-- -172
x"fe990",-- -359
x"fe710",-- -399
x"fe1c0",-- -484
x"fd7c0",-- -644
x"fd850",-- -635
x"fd5d0",-- -675
x"fd200",-- -736
x"fd360",-- -714
x"fca80",-- -856
x"fce10",-- -799
x"fcfa0",-- -774
x"fca20",-- -862
x"fd1b0",-- -741
x"fd4c0",-- -692
x"fd1d0",-- -739
x"fcfa0",-- -774
x"fcff0",-- -769
x"fd4c0",-- -692
x"fd020",-- -766
x"fcbc0",-- -836
x"fd020",-- -766
x"fccb0",-- -821
x"fd100",-- -752
x"fd440",-- -700
x"fd400",-- -704
x"fd720",-- -654
x"fda10",-- -607
x"fd880",-- -632
x"fd850",-- -635
x"fd5b0",-- -677
x"fd790",-- -647
x"fdab0",-- -597
x"fd5d0",-- -675
x"fdb80",-- -584
x"fe140",-- -492
x"fe730",-- -397
x"fea80",-- -344
x"fef00",-- -272
x"fecd0",-- -307
x"fecf0",-- -305
x"ff380",-- -200
x"ff7b0",-- -133
x"ffdd0",-- -35
x"fffe0",-- -2
x"00320",-- 50
x"00570",-- 87
x"00700",-- 112
x"00c00",-- 192
x"00de0",-- 222
x"00d90",-- 217
x"00e60",-- 230
x"01180",-- 280
x"013d0",-- 317
x"016c0",-- 364
x"01b70",-- 439
x"01b70",-- 439
x"01a90",-- 425
x"01d00",-- 464
x"01b70",-- 439
x"01c20",-- 450
x"01e20",-- 482
x"01c10",-- 449
x"01d30",-- 467
x"01e50",-- 485
x"01a10",-- 417
x"01950",-- 405
x"01740",-- 372
x"019e0",-- 414
x"01990",-- 409
x"016d0",-- 365
x"01a60",-- 422
x"017c0",-- 380
x"01510",-- 337
x"01220",-- 290
x"013f0",-- 319
x"01630",-- 355
x"01470",-- 327
x"01630",-- 355
x"01990",-- 409
x"01d10",-- 465
x"01dd0",-- 477
x"020f0",-- 527
x"022b0",-- 555
x"024b0",-- 587
x"02460",-- 582
x"02640",-- 612
x"02a20",-- 674
x"029d0",-- 669
x"02f40",-- 756
x"034a0",-- 842
x"03420",-- 834
x"03990",-- 921
x"03f80",-- 1016
x"04490",-- 1097
x"04980",-- 1176
x"04c70",-- 1223
x"048f0",-- 1167
x"04320",-- 1074
x"03b70",-- 951
x"03a30",-- 931
x"03090",-- 777
x"02170",-- 535
x"01560",-- 342
x"00c00",-- 192
x"005a0",-- 90
x"ffee0",-- -18
x"ffb20",-- -78
x"ff530",-- -173
x"ff020",-- -254
x"fe890",-- -375
x"fe300",-- -464
x"fe050",-- -507
x"fd950",-- -619
x"fce90",-- -791
x"fc430",-- -957
x"fbc90",-- -1079
x"fb970",-- -1129
x"fb970",-- -1129
x"fb570",-- -1193
x"fb1f0",-- -1249
x"fb600",-- -1184
x"fbb30",-- -1101
x"fc0d0",-- -1011
x"fc5f0",-- -929
x"fcb10",-- -847
x"fce60",-- -794
x"fd020",-- -766
x"fcfd0",-- -771
x"fd2f0",-- -721
x"fd4f0",-- -689
x"fd3a0",-- -710
x"fd2f0",-- -721
x"fd1b0",-- -741
x"fd4e0",-- -690
x"fd6c0",-- -660
x"fd800",-- -640
x"fd970",-- -617
x"fda80",-- -600
x"fd940",-- -620
x"fd6f0",-- -657
x"fd4e0",-- -690
x"fd630",-- -669
x"fd710",-- -655
x"fd2a0",-- -726
x"fd200",-- -736
x"fd440",-- -700
x"fd8f0",-- -625
x"fdd10",-- -559
x"fdd30",-- -557
x"fe160",-- -490
x"fe530",-- -429
x"fea20",-- -350
x"fe9b0",-- -357
x"fe840",-- -380
x"fec10",-- -319
x"ff0c0",-- -244
x"ff1c0",-- -228
x"ff2c0",-- -212
x"ff7b0",-- -133
x"ffab0",-- -85
x"ffc20",-- -62
x"ff4a0",-- -182
x"ffbc0",-- -68
x"00390",-- 57
x"fffd0",-- -3
x"00120",-- 18
x"003e0",-- 62
x"00430",-- 67
x"00940",-- 148
x"00840",-- 132
x"00670",-- 103
x"00b20",-- 178
x"00a70",-- 167
x"006c0",-- 108
x"007a0",-- 122
x"00dc0",-- 220
x"00e10",-- 225
x"00a80",-- 168
x"007d0",-- 125
x"007d0",-- 125
x"00800",-- 128
x"00b10",-- 177
x"00eb0",-- 235
x"00f90",-- 249
x"01240",-- 292
x"01310",-- 305
x"01180",-- 280
x"01450",-- 325
x"01600",-- 352
x"01590",-- 345
x"01680",-- 360
x"01a90",-- 425
x"01c60",-- 454
x"01d10",-- 465
x"022b0",-- 555
x"02890",-- 649
x"02c00",-- 704
x"031f0",-- 799
x"03180",-- 792
x"03850",-- 901
x"03da0",-- 986
x"041e0",-- 1054
x"04b80",-- 1208
x"05360",-- 1334
x"05b80",-- 1464
x"06460",-- 1606
x"06fc0",-- 1788
x"07c60",-- 1990
x"08a20",-- 2210
x"09bf0",-- 2495
x"09f80",-- 2552
x"09470",-- 2375
x"08680",-- 2152
x"07f80",-- 2040
x"07150",-- 1813
x"056a0",-- 1386
x"03880",-- 904
x"01970",-- 407
x"00480",-- 72
x"fefc0",-- -260
x"fde70",-- -537
x"fd2c0",-- -724
x"fcb40",-- -844
x"fc020",-- -1022
x"fb6f0",-- -1169
x"fb770",-- -1161
x"fb600",-- -1184
x"fac30",-- -1341
x"f9e90",-- -1559
x"f91d0",-- -1763
x"f8da0",-- -1830
x"f9090",-- -1783
x"f9040",-- -1788
x"f91a0",-- -1766
x"f9ab0",-- -1621
x"fab20",-- -1358
x"fb9c0",-- -1124
x"fcaf0",-- -849
x"fda60",-- -602
x"fe520",-- -430
x"fe9b0",-- -357
x"feb60",-- -330
x"ff2e0",-- -210
x"ff5d0",-- -163
x"ff290",-- -215
x"fe9b0",-- -357
x"fe460",-- -442
x"fe580",-- -424
x"fe750",-- -395
x"fe3c0",-- -452
x"fe140",-- -492
x"fde70",-- -537
x"fdbd0",-- -579
x"fdc10",-- -575
x"fd9a0",-- -614
x"fd810",-- -639
x"fd3a0",-- -710
x"fcd70",-- -809
x"fcaa0",-- -854
x"fcc30",-- -829
x"fcfd0",-- -771
x"fd1a0",-- -742
x"fcff0",-- -769
x"fd530",-- -685
x"fd240",-- -732
x"fd110",-- -751
x"fdc10",-- -575
x"fe0d0",-- -499
x"fe440",-- -444
x"fe490",-- -439
x"fe9e0",-- -354
x"fef80",-- -264
x"fee90",-- -279
x"ff470",-- -185
x"ff4e0",-- -178
x"ff970",-- -105
x"ff8a0",-- -118
x"ff4f0",-- -177
x"ffc40",-- -60
x"00000",-- 0
x"ffe20",-- -30
x"ff540",-- -172
x"ff720",-- -142
x"ffea0",-- -22
x"fff60",-- -10
x"00280",-- 40
x"001e0",-- 30
x"00530",-- 83
x"00700",-- 112
x"00750",-- 117
x"00120",-- 18
x"00210",-- 33
x"ffec0",-- -20
x"fee40",-- -284
x"ff6a0",-- -150
x"ff790",-- -135
x"ffc40",-- -60
x"006e0",-- 110
x"00a70",-- 167
x"00ca0",-- 202
x"011f0",-- 287
x"01880",-- 392
x"017b0",-- 379
x"018b0",-- 395
x"02430",-- 579
x"02320",-- 562
x"02a70",-- 679
x"02cc0",-- 716
x"03290",-- 809
x"03e00",-- 992
x"04000",-- 1024
x"04bb0",-- 1211
x"05630",-- 1379
x"06280",-- 1576
x"06b10",-- 1713
x"073b0",-- 1851
x"084b0",-- 2123
x"09170",-- 2327
x"0a390",-- 2617
x"0b860",-- 2950
x"0ce60",-- 3302
x"0ed10",-- 3793
x"10550",-- 4181
x"11bc0",-- 4540
x"12390",-- 4665
x"11fa0",-- 4602
x"11040",-- 4356
x"0f650",-- 3941
x"0d150",-- 3349
x"09b70",-- 2487
x"05ae0",-- 1454
x"019e0",-- 414
x"fdf80",-- -520
x"fa7a0",-- -1414
x"f7540",-- -2220
x"f4c30",-- -2877
x"f2930",-- -3437
x"f12c0",-- -3796
x"f08e0",-- -3954
x"f0730",-- -3981
x"f0a50",-- -3931
x"f0d70",-- -3881
x"f1090",-- -3831
x"f1980",-- -3688
x"f29b0",-- -3429
x"f3d10",-- -3119
x"f4dc0",-- -2852
x"f66c0",-- -2452
x"f8570",-- -1961
x"fab20",-- -1358
x"fd670",-- -665
x"00200",-- 32
x"02710",-- 625
x"049e0",-- 1182
x"06610",-- 1633
x"07970",-- 1943
x"08640",-- 2148
x"08520",-- 2130
x"07770",-- 1911
x"06210",-- 1569
x"04930",-- 1171
x"02c30",-- 707
x"00f50",-- 245
x"fefa0",-- -262
x"fd090",-- -759
x"fb590",-- -1191
x"fa0d0",-- -1523
x"f8e80",-- -1816
x"f7f40",-- -2060
x"f7380",-- -2248
x"f68f0",-- -2417
x"f6250",-- -2523
x"f61e0",-- -2530
x"f6280",-- -2520
x"f67d0",-- -2435
x"f6c00",-- -2368
x"f77c0",-- -2180
x"f8000",-- -2048
x"f8ad0",-- -1875
x"f9a10",-- -1631
x"faa80",-- -1368
x"fc1c0",-- -996
x"fd3f0",-- -705
x"feb20",-- -334
x"004b0",-- 75
x"01fd0",-- 509
x"03560",-- 854
x"04110",-- 1041
x"04cc0",-- 1228
x"05040",-- 1284
x"04a70",-- 1191
x"04170",-- 1047
x"033f0",-- 831
x"02800",-- 640
x"01400",-- 320
x"00250",-- 37
x"ff540",-- -172
x"fede0",-- -290
x"fe690",-- -407
x"fdda0",-- -550
x"fda90",-- -599
x"fd990",-- -615
x"fda10",-- -607
x"fd830",-- -637
x"fd680",-- -664
x"fd400",-- -704
x"fcf70",-- -777
x"fcb70",-- -841
x"fca20",-- -862
x"fd090",-- -759
x"fd650",-- -667
x"fdfb0",-- -517
x"fede0",-- -290
x"00320",-- 50
x"01bd0",-- 445
x"03100",-- 784
x"04390",-- 1081
x"05350",-- 1333
x"063a0",-- 1594
x"06d20",-- 1746
x"07220",-- 1826
x"074f0",-- 1871
x"07740",-- 1908
x"079c0",-- 1948
x"07e70",-- 2023
x"088c0",-- 2188
x"091a0",-- 2330
x"09e40",-- 2532
x"0ac80",-- 2760
x"0c1b0",-- 3099
x"0dec0",-- 3564
x"0fe70",-- 4071
x"12270",-- 4647
x"14000",-- 5120
x"15aa0",-- 5546
x"17100",-- 5904
x"188b0",-- 6283
x"18d20",-- 6354
x"17d50",-- 6101
x"155b0",-- 5467
x"12130",-- 4627
x"0dbd0",-- 3517
x"08ac0",-- 2220
x"02c80",-- 712
x"fcc30",-- -829
x"f72a0",-- -2262
x"f1d10",-- -3631
x"edce0",-- -4658
x"ea510",-- -5551
x"e82e0",-- -6098
x"e6500",-- -6576
x"e5510",-- -6831
x"e60b0",-- -6645
x"e76d0",-- -6291
x"e9700",-- -5776
x"eb110",-- -5359
x"ed630",-- -4765
x"eff90",-- -4103
x"f2af0",-- -3409
x"f5ca0",-- -2614
x"f8cf0",-- -1841
x"fbf30",-- -1037
x"ff9c0",-- -100
x"03440",-- 836
x"06cc0",-- 1740
x"0a460",-- 2630
x"0d210",-- 3361
x"0ee60",-- 3814
x"0fcb0",-- 4043
x"0fe20",-- 4066
x"0eed0",-- 3821
x"0ce00",-- 3296
x"09b50",-- 2485
x"062d0",-- 1581
x"028e0",-- 654
x"fec50",-- -315
x"fab90",-- -1351
x"f7160",-- -2282
x"f4070",-- -3065
x"f1c50",-- -3643
x"efc70",-- -4153
x"ee8e0",-- -4466
x"eddd0",-- -4643
x"ed9a0",-- -4710
x"eda10",-- -4703
x"ee260",-- -4570
x"ef2a0",-- -4310
x"f06b0",-- -3989
x"f2100",-- -3568
x"f3b30",-- -3149
x"f6030",-- -2557
x"f8b20",-- -1870
x"fbc70",-- -1081
x"feb40",-- -332
x"025d0",-- 605
x"05030",-- 1283
x"07dd0",-- 2013
x"0a320",-- 2610
x"0c370",-- 3127
x"0d970",-- 3479
x"0de40",-- 3556
x"0ccd0",-- 3277
x"0b560",-- 2902
x"09f10",-- 2545
x"07260",-- 1830
x"04140",-- 1044
x"00cb0",-- 203
x"fdfd0",-- -515
x"fb480",-- -1208
x"f92f0",-- -1745
x"f73e0",-- -2242
x"f6300",-- -2512
x"f5c00",-- -2624
x"f54a0",-- -2742
x"f5570",-- -2729
x"f65a0",-- -2470
x"f70c0",-- -2292
x"f7b50",-- -2123
x"f8410",-- -1983
x"f95e0",-- -1698
x"fa870",-- -1401
x"fbc60",-- -1082
x"fcf70",-- -777
x"fe200",-- -480
x"003f0",-- 63
x"028a0",-- 650
x"04980",-- 1176
x"06be0",-- 1726
x"08d70",-- 2263
x"0ab40",-- 2740
x"0bd50",-- 3029
x"0ce00",-- 3296
x"0d470",-- 3399
x"0d470",-- 3399
x"0c960",-- 3222
x"0b7e0",-- 2942
x"0a6e0",-- 2670
x"09e00",-- 2528
x"08f50",-- 2293
x"08430",-- 2115
x"08720",-- 2162
x"09770",-- 2423
x"0adb0",-- 2779
x"0d240",-- 3364
x"10570",-- 4183
x"13820",-- 4994
x"16500",-- 5712
x"182d0",-- 6189
x"1a070",-- 6663
x"1b5f0",-- 7007
x"1b740",-- 7028
x"18860",-- 6278
x"165a0",-- 5722
x"13990",-- 5017
x"0d4c0",-- 3404
x"06610",-- 1633
x"fe3a0",-- -454
x"f69b0",-- -2405
x"effc0",-- -4100
x"e9bd0",-- -5699
x"e50e0",-- -6898
x"e26f0",-- -7569
x"e25d0",-- -7587
x"e26a0",-- -7574
x"e3480",-- -7352
x"e5980",-- -6760
x"e8410",-- -6079
x"eaf20",-- -5390
x"ed1b0",-- -4837
x"ef610",-- -4255
x"f27f0",-- -3457
x"f62b0",-- -2517
x"f9790",-- -1671
x"fd360",-- -714
x"01900",-- 400
x"05b30",-- 1459
x"09b80",-- 2488
x"0d7b0",-- 3451
x"10cc0",-- 4300
x"132b0",-- 4907
x"13bc0",-- 5052
x"12cc0",-- 4812
x"10e80",-- 4328
x"0db70",-- 3511
x"09330",-- 2355
x"03920",-- 914
x"fd630",-- -669
x"f8200",-- -2016
x"f3390",-- -3271
x"eed90",-- -4391
x"eb630",-- -5277
x"e97e0",-- -5762
x"e8c10",-- -5951
x"e8ed0",-- -5907
x"e9950",-- -5739
x"eb270",-- -5337
x"ed020",-- -4862
x"ef220",-- -4318
x"f0fa0",-- -3846
x"f2e40",-- -3356
x"f4e60",-- -2842
x"f7980",-- -2152
x"fa500",-- -1456
x"fce90",-- -791
x"ffc90",-- -55
x"039e0",-- 926
x"07c90",-- 1993
x"0b6f0",-- 2927
x"0eb60",-- 3766
x"11560",-- 4438
x"13960",-- 5014
x"146b0",-- 5227
x"13770",-- 4983
x"11900",-- 4496
x"0e8b0",-- 3723
x"09d50",-- 2517
x"04c70",-- 1223
x"ffd00",-- -48
x"fb5b0",-- -1189
x"f6a20",-- -2398
x"f2dc0",-- -3364
x"f09d0",-- -3939
x"f0120",-- -4078
x"f0640",-- -3996
x"f0f50",-- -3851
x"f26e0",-- -3474
x"f4c10",-- -2879
x"f7150",-- -2283
x"f8b70",-- -1865
x"f9cc0",-- -1588
x"faf30",-- -1293
x"fbfd0",-- -1027
x"fccd0",-- -819
x"fd800",-- -640
x"fe960",-- -362
x"004b0",-- 75
x"02320",-- 562
x"041e0",-- 1054
x"06930",-- 1683
x"09220",-- 2338
x"0b2b0",-- 2859
x"0c570",-- 3159
x"0d4f0",-- 3407
x"0dc90",-- 3529
x"0d740",-- 3444
x"0c190",-- 3097
x"0a260",-- 2598
x"08840",-- 2180
x"06d70",-- 1751
x"05210",-- 1313
x"03a90",-- 937
x"032c0",-- 812
x"039c0",-- 924
x"04ca0",-- 1226
x"06cc0",-- 1740
x"09b00",-- 2480
x"0d1f0",-- 3359
x"11420",-- 4418
x"14e00",-- 5344
x"185a0",-- 6234
x"1b230",-- 6947
x"1d0f0",-- 7439
x"1e230",-- 7715
x"1d560",-- 7510
x"1b9b0",-- 7067
x"17730",-- 6003
x"13150",-- 4885
x"0d270",-- 3367
x"06730",-- 1651
x"ff670",-- -153
x"f8570",-- -1961
x"f2370",-- -3529
x"ec420",-- -5054
x"e80f0",-- -6129
x"e43c0",-- -7108
x"e2640",-- -7580
x"e1570",-- -7849
x"e1540",-- -7852
x"e2230",-- -7645
x"e3e00",-- -7200
x"e6790",-- -6535
x"e91f0",-- -5857
x"eca50",-- -4955
x"f0760",-- -3978
x"f5150",-- -2795
x"f99f0",-- -1633
x"fe890",-- -375
x"03630",-- 867
x"083c0",-- 2108
x"0c9b0",-- 3227
x"10070",-- 4103
x"129d0",-- 4765
x"14250",-- 5157
x"14690",-- 5225
x"13150",-- 4885
x"10770",-- 4215
x"0cd10",-- 3281
x"08690",-- 2153
x"03650",-- 869
x"fe170",-- -489
x"f8cb0",-- -1845
x"f40c0",-- -3060
x"efe00",-- -4128
x"ec8e0",-- -4978
x"ea380",-- -5576
x"e8b00",-- -5968
x"e7fe0",-- -6146
x"e8030",-- -6141
x"e8e90",-- -5911
x"ea910",-- -5487
x"ec1a0",-- -5094
x"ee240",-- -4572
x"f09b0",-- -3941
x"f3ec0",-- -3092
x"f7520",-- -2222
x"fae10",-- -1311
x"fea30",-- -349
x"02ea0",-- 746
x"07620",-- 1890
x"0b7e0",-- 2942
x"0f4f0",-- 3919
x"125f0",-- 4703
x"14b90",-- 5305
x"15c30",-- 5571
x"15c10",-- 5569
x"14720",-- 5234
x"12390",-- 4665
x"0eaa0",-- 3754
x"0a110",-- 2577
x"051f0",-- 1311
x"00570",-- 87
x"fbcb0",-- -1077
x"f7250",-- -2267
x"f36b0",-- -3221
x"f0cd0",-- -3891
x"efa10",-- -4191
x"ef2e0",-- -4306
x"ef2e0",-- -4306
x"eff90",-- -4103
x"f1c00",-- -3648
x"f3d60",-- -3114
x"f5c00",-- -2624
x"f7d00",-- -2096
x"f9970",-- -1641
x"fb420",-- -1214
x"fcf50",-- -779
x"febb0",-- -325
x"00890",-- 137
x"024b0",-- 587
x"04230",-- 1059
x"061b0",-- 1563
x"08640",-- 2148
x"0a7c0",-- 2684
x"0bee0",-- 3054
x"0ca50",-- 3237
x"0d270",-- 3367
x"0d2b0",-- 3371
x"0c7d0",-- 3197
x"0b010",-- 2817
x"09270",-- 2343
x"06ed0",-- 1773
x"05240",-- 1316
x"03210",-- 801
x"01ba0",-- 442
x"00710",-- 113
x"00350",-- 53
x"00800",-- 128
x"01f10",-- 497
x"04170",-- 1047
x"068c0",-- 1676
x"0a0c0",-- 2572
x"0dad0",-- 3501
x"12040",-- 4612
x"15350",-- 5429
x"18840",-- 6276
x"1ac80",-- 6856
x"1cef0",-- 7407
x"1e140",-- 7700
x"1d920",-- 7570
x"1c2d0",-- 7213
x"18e10",-- 6369
x"14ea0",-- 5354
x"0fd50",-- 4053
x"0a300",-- 2608
x"03360",-- 822
x"fbba0",-- -1094
x"f5200",-- -2784
x"eec00",-- -4416
x"e9bf0",-- -5697
x"e4b40",-- -6988
x"e1280",-- -7896
x"ded70",-- -8489
x"de4b0",-- -8629
x"dee60",-- -8474
x"e04c0",-- -8116
x"e2e10",-- -7455
x"e6150",-- -6635
x"eaa60",-- -5466
x"ef740",-- -4236
x"f4d50",-- -2859
x"f9d30",-- -1581
x"fee80",-- -280
x"03f60",-- 1014
x"088b0",-- 2187
x"0ca70",-- 3239
x"0f800",-- 3968
x"118b0",-- 4491
x"125a0",-- 4698
x"12de0",-- 4830
x"11df0",-- 4575
x"0fe20",-- 4066
x"0cd70",-- 3287
x"09220",-- 2338
x"054c0",-- 1356
x"01090",-- 265
x"fca20",-- -862
x"f7d60",-- -2090
x"f3cf0",-- -3121
x"efea0",-- -4118
x"ecdc0",-- -4900
x"ea260",-- -5594
x"e8210",-- -6111
x"e6b90",-- -6471
x"e66f0",-- -6545
x"e76f0",-- -6289
x"e91a0",-- -5862
x"eb5c0",-- -5284
x"ee700",-- -4496
x"f2460",-- -3514
x"f6de0",-- -2338
x"fbc90",-- -1079
x"00750",-- 117
x"04eb0",-- 1259
x"093d0",-- 2365
x"0d6d0",-- 3437
x"10a20",-- 4258
x"13130",-- 4883
x"13f00",-- 5104
x"14250",-- 5157
x"13dc0",-- 5084
x"12860",-- 4742
x"10430",-- 4163
x"0cc50",-- 3269
x"08f90",-- 2297
x"05400",-- 1344
x"019e0",-- 414
x"fd970",-- -617
x"f9420",-- -1726
x"f6160",-- -2538
x"f3750",-- -3211
x"f1c20",-- -3646
x"f0460",-- -4026
x"ef890",-- -4215
x"ef790",-- -4231
x"f06b0",-- -3989
x"f18d0",-- -3699
x"f3420",-- -3262
x"f5750",-- -2699
x"f7600",-- -2208
x"f99c0",-- -1636
x"fc0d0",-- -1011
x"fef20",-- -270
x"01770",-- 375
x"038f0",-- 911
x"057c0",-- 1404
x"078d0",-- 1933
x"09cb0",-- 2507
x"0b060",-- 2822
x"0b810",-- 2945
x"0b940",-- 2964
x"0bd00",-- 3024
x"0b680",-- 2920
x"0a200",-- 2592
x"08720",-- 2162
x"06af0",-- 1711
x"05270",-- 1319
x"038d0",-- 909
x"01df0",-- 479
x"00840",-- 132
x"ffd30",-- -45
x"ff6f0",-- -145
x"ff990",-- -103
x"00840",-- 132
x"02120",-- 530
x"03e90",-- 1001
x"06670",-- 1639
x"09720",-- 2418
x"0cf50",-- 3317
x"10f20",-- 4338
x"141e0",-- 5150
x"16d70",-- 5847
x"196f0",-- 6511
x"1c070",-- 7175
x"1dec0",-- 7660
x"1da00",-- 7584
x"1ca70",-- 7335
x"19c30",-- 6595
x"17460",-- 5958
x"12c30",-- 4803
x"0caf0",-- 3247
x"055d0",-- 1373
x"fe000",-- -512
x"f7860",-- -2170
x"f04b0",-- -4021
x"ea870",-- -5497
x"e4080",-- -7160
x"e0650",-- -8091
x"ddbb0",-- -8773
x"dcd00",-- -9008
x"dcc80",-- -9016
x"de300",-- -8656
x"e11e0",-- -7906
x"e4880",-- -7032
x"e9d90",-- -5671
x"eed00",-- -4400
x"f46e0",-- -2962
x"f98d0",-- -1651
x"feaf0",-- -337
x"03d50",-- 981
x"08730",-- 2163
x"0bfd0",-- 3069
x"0e070",-- 3591
x"0ffd0",-- 4093
x"11330",-- 4403
x"11da0",-- 4570
x"10cc0",-- 4300
x"0ed90",-- 3801
x"0ca20",-- 3234
x"0a480",-- 2632
x"07770",-- 1911
x"03970",-- 919
x"ff8d0",-- -115
x"fbb70",-- -1097
x"f8300",-- -2000
x"f46b0",-- -2965
x"f1040",-- -3836
x"edf10",-- -4623
x"eb630",-- -5277
x"e9d40",-- -5676
x"e8e10",-- -5919
x"e8f30",-- -5901
x"e9c50",-- -5691
x"eb750",-- -5259
x"edb00",-- -4688
x"f1160",-- -3818
x"f5020",-- -2814
x"f90c0",-- -1780
x"fd4a0",-- -694
x"01400",-- 320
x"059c0",-- 1436
x"09740",-- 2420
x"0ce60",-- 3302
x"0eea0",-- 3818
x"10cf0",-- 4303
x"120a0",-- 4618
x"12820",-- 4738
x"12340",-- 4660
x"108e0",-- 4238
x"0ee60",-- 3814
x"0c820",-- 3202
x"0a000",-- 2560
x"06cc0",-- 1740
x"02480",-- 584
x"ff1d0",-- -227
x"fb400",-- -1216
x"f8a20",-- -1886
x"f4e90",-- -2839
x"f23f0",-- -3521
x"f05d0",-- -4003
x"ef330",-- -4301
x"ef4d0",-- -4275
x"ee700",-- -4496
x"efe80",-- -4120
x"f1090",-- -3831
x"f38d0",-- -3187
x"f5c20",-- -2622
x"f88c0",-- -1908
x"fb8b0",-- -1141
x"fe0f0",-- -497
x"010b0",-- 267
x"03580",-- 856
x"05f30",-- 1523
x"07b50",-- 1973
x"08b60",-- 2230
x"09a40",-- 2468
x"0a080",-- 2568
x"0a590",-- 2649
x"09590",-- 2393
x"08500",-- 2128
x"07090",-- 1801
x"06300",-- 1584
x"04e80",-- 1256
x"037b0",-- 891
x"02230",-- 547
x"017b0",-- 379
x"01030",-- 259
x"00a30",-- 163
x"00520",-- 82
x"00b10",-- 177
x"01650",-- 357
x"02390",-- 569
x"03c40",-- 964
x"05790",-- 1401
x"07d60",-- 2006
x"0a0d0",-- 2573
x"0cdc0",-- 3292
x"10070",-- 4103
x"13080",-- 4872
x"15c30",-- 5571
x"17d20",-- 6098
x"1a810",-- 6785
x"1c4d0",-- 7245
x"1caa0",-- 7338
x"1c2c0",-- 7212
x"1a050",-- 6661
x"17d80",-- 6104
x"13740",-- 4980
x"0ebb0",-- 3771
x"07c90",-- 1993
x"01290",-- 297
x"faa30",-- -1373
x"f39d0",-- -3171
x"eda10",-- -4703
x"e7570",-- -6313
x"e34c0",-- -7348
x"df750",-- -8331
x"de3d0",-- -8643
x"dd720",-- -8846
x"de240",-- -8668
x"e0760",-- -8074
x"e3790",-- -7303
x"e7f60",-- -6154
x"eca30",-- -4957
x"f22a0",-- -3542
x"f6fa0",-- -2310
x"fc550",-- -939
x"01580",-- 344
x"05c10",-- 1473
x"094f0",-- 2383
x"0bec0",-- 3052
x"0dcc0",-- 3532
x"0f1a0",-- 3866
x"0fa40",-- 4004
x"0f0e0",-- 3854
x"0dd10",-- 3537
x"0c190",-- 3097
x"0a3c0",-- 2620
x"07d00",-- 2000
x"05310",-- 1329
x"02120",-- 530
x"ff220",-- -222
x"fc490",-- -951
x"f98d0",-- -1651
x"f6b10",-- -2383
x"f3fb0",-- -3077
x"f1ec0",-- -3604
x"f00b0",-- -4085
x"eebe0",-- -4418
x"edec0",-- -4628
x"ed860",-- -4730
x"edcf0",-- -4657
x"eeb60",-- -4426
x"f0520",-- -4014
x"f2870",-- -3449
x"f5220",-- -2782
x"f8000",-- -2048
x"fb570",-- -1193
x"fecb0",-- -309
x"02320",-- 562
x"05590",-- 1369
x"085f0",-- 2143
x"0ae60",-- 2790
x"0cf90",-- 3321
x"0e810",-- 3713
x"0f7e0",-- 3966
x"0fee0",-- 4078
x"0f9f0",-- 3999
x"0ecf0",-- 3791
x"0d1a0",-- 3354
x"0b240",-- 2852
x"08f90",-- 2297
x"05bf0",-- 1471
x"02480",-- 584
x"fee80",-- -280
x"fb9e0",-- -1122
x"f8b40",-- -1868
x"f5330",-- -2765
x"f2c80",-- -3384
x"f0890",-- -3959
x"efca0",-- -4150
x"ef1d0",-- -4323
x"eeb40",-- -4428
x"efe70",-- -4121
x"f1560",-- -3754
x"f3bd0",-- -3139
x"f5e90",-- -2583
x"f8cd0",-- -1843
x"fbc90",-- -1079
x"fea20",-- -350
x"01710",-- 369
x"03620",-- 866
x"05800",-- 1408
x"06ef0",-- 1775
x"07c10",-- 1985
x"08210",-- 2081
x"080f0",-- 2063
x"08210",-- 2081
x"07180",-- 1816
x"067d0",-- 1661
x"058b0",-- 1419
x"04e10",-- 1249
x"04340",-- 1076
x"03330",-- 819
x"02af0",-- 687
x"02750",-- 629
x"028c0",-- 652
x"024e0",-- 590
x"02140",-- 532
x"02930",-- 659
x"03210",-- 801
x"039f0",-- 927
x"04750",-- 1141
x"05380",-- 1336
x"07010",-- 1793
x"08840",-- 2180
x"0abd0",-- 2749
x"0cd70",-- 3287
x"0f470",-- 3911
x"121b0",-- 4635
x"14410",-- 5185
x"16be0",-- 5822
x"185a0",-- 6234
x"19850",-- 6533
x"19c90",-- 6601
x"18c70",-- 6343
x"17780",-- 6008
x"14610",-- 5217
x"109b0",-- 4251
x"0b830",-- 2947
x"05a30",-- 1443
x"00250",-- 37
x"f96a0",-- -1686
x"f3ac0",-- -3156
x"ed1b0",-- -4837
x"e8780",-- -6024
x"e45d0",-- -7075
x"e1610",-- -7839
x"df980",-- -8296
x"de8c0",-- -8564
x"dfec0",-- -8212
x"e1b60",-- -7754
x"e52f0",-- -6865
x"e8d00",-- -5936
x"ed8e0",-- -4722
x"f2b60",-- -3402
x"f7e50",-- -2075
x"fd010",-- -767
x"017e0",-- 382
x"05b50",-- 1461
x"09040",-- 2308
x"0bb20",-- 2994
x"0d4c0",-- 3404
x"0e430",-- 3651
x"0e3b0",-- 3643
x"0da80",-- 3496
x"0c630",-- 3171
x"0abd0",-- 2749
x"08c30",-- 2243
x"06640",-- 1636
x"04070",-- 1031
x"017b0",-- 379
x"ff740",-- -140
x"fd1b0",-- -741
x"fafd0",-- -1283
x"f8eb0",-- -1813
x"f7590",-- -2215
x"f6110",-- -2543
x"f4c10",-- -2879
x"f3c40",-- -3132
x"f2c10",-- -3391
x"f27d0",-- -3459
x"f2500",-- -3504
x"f27a0",-- -3462
x"f2de0",-- -3362
x"f3a60",-- -3162
x"f5220",-- -2782
x"f6b60",-- -2378
x"f8f20",-- -1806
x"fb310",-- -1231
x"fdda0",-- -550
x"00a80",-- 168
x"03ab0",-- 939
x"06930",-- 1683
x"08f50",-- 2293
x"0b440",-- 2884
x"0cf90",-- 3321
x"0e5c0",-- 3676
x"0f090",-- 3849
x"0ef40",-- 3828
x"0e430",-- 3651
x"0cc50",-- 3269
x"0ae10",-- 2785
x"086e0",-- 2158
x"05590",-- 1369
x"01e00",-- 480
x"fe690",-- -407
x"fb110",-- -1263
x"f8140",-- -2028
x"f5010",-- -2815
x"f2bc0",-- -3396
x"f0cf0",-- -3889
x"f00a0",-- -4086
x"efd40",-- -4140
x"eff10",-- -4111
x"f0fc0",-- -3844
x"f2570",-- -3497
x"f4930",-- -2925
x"f6af0",-- -2385
x"f9360",-- -1738
x"fb7b0",-- -1157
x"fe070",-- -505
x"00550",-- 85
x"02480",-- 584
x"03c60",-- 966
x"04f50",-- 1269
x"05bc0",-- 1468
x"06300",-- 1584
x"06440",-- 1604
x"06230",-- 1571
x"05b50",-- 1461
x"051d0",-- 1309
x"04b40",-- 1204
x"040a0",-- 1034
x"03bf0",-- 959
x"03310",-- 817
x"02f20",-- 754
x"02cd0",-- 717
x"03170",-- 791
x"03450",-- 837
x"03650",-- 869
x"03c90",-- 969
x"04550",-- 1109
x"04fe0",-- 1278
x"05a60",-- 1446
x"06620",-- 1634
x"07470",-- 1863
x"08a50",-- 2213
x"0a300",-- 2608
x"0c1d0",-- 3101
x"0db00",-- 3504
x"0fee0",-- 4078
x"119f0",-- 4511
x"13e20",-- 5090
x"15850",-- 5509
x"16900",-- 5776
x"171c0",-- 5916
x"16720",-- 5746
x"163b0",-- 5691
x"13ad0",-- 5037
x"11580",-- 4440
x"0ce10",-- 3297
x"08960",-- 2198
x"03fb0",-- 1019
x"fe710",-- -399
x"f92f0",-- -1745
x"f2ee0",-- -3346
x"ee910",-- -4463
x"ea000",-- -5632
x"e6a80",-- -6488
x"e3880",-- -7288
x"e1ba0",-- -7750
x"e1810",-- -7807
x"e1fe0",-- -7682
x"e3f40",-- -7180
x"e61e0",-- -6626
x"e9db0",-- -5669
x"ede30",-- -4637
x"f2990",-- -3431
x"f7590",-- -2215
x"fc190",-- -999
x"00990",-- 153
x"047b0",-- 1147
x"08200",-- 2080
x"0aca0",-- 2762
x"0cef0",-- 3311
x"0dda0",-- 3546
x"0e360",-- 3638
x"0da60",-- 3494
x"0cc80",-- 3272
x"0b440",-- 2884
x"08fe0",-- 2302
x"06af0",-- 1711
x"042d0",-- 1069
x"02210",-- 545
x"ffc20",-- -62
x"fd8f0",-- -625
x"fb9a0",-- -1126
x"f9f60",-- -1546
x"f8f70",-- -1801
x"f7920",-- -2158
x"f6e10",-- -2335
x"f5e20",-- -2590
x"f5bd0",-- -2627
x"f58e0",-- -2674
x"f5520",-- -2734
x"f59d0",-- -2659
x"f5930",-- -2669
x"f6700",-- -2448
x"f6fa0",-- -2310
x"f83e0",-- -1986
x"f9830",-- -1661
x"fb110",-- -1263
x"fced0",-- -787
x"fede0",-- -290
x"01350",-- 309
x"03490",-- 841
x"055b0",-- 1371
x"07420",-- 1858
x"09290",-- 2345
x"0aae0",-- 2734
x"0ba80",-- 2984
x"0bdf0",-- 3039
x"0bdf0",-- 3039
x"0b880",-- 2952
x"0ab30",-- 2739
x"09420",-- 2370
x"06be0",-- 1726
x"04f50",-- 1269
x"022f0",-- 559
x"ffd00",-- -48
x"fcaf0",-- -849
x"f9c20",-- -1598
x"f7c10",-- -2111
x"f5110",-- -2799
x"f3e80",-- -3096
x"f1a90",-- -3671
x"f1560",-- -3754
x"f0e30",-- -3869
x"f0f30",-- -3853
x"f1f40",-- -3596
x"f2a00",-- -3424
x"f4b20",-- -2894
x"f61e0",-- -2530
x"f86e0",-- -1938
x"fa960",-- -1386
x"fced0",-- -787
x"ff4c0",-- -180
x"011c0",-- 284
x"03010",-- 769
x"049d0",-- 1181
x"05fe0",-- 1534
x"06cd0",-- 1741
x"070b0",-- 1803
x"07540",-- 1876
x"07380",-- 1848
x"06c80",-- 1736
x"06050",-- 1541
x"05240",-- 1316
x"046c0",-- 1132
x"03e50",-- 997
x"032c0",-- 812
x"02c00",-- 704
x"026e0",-- 622
x"02940",-- 660
x"02cc0",-- 716
x"03260",-- 806
x"03e40",-- 996
x"04890",-- 1161
x"05b50",-- 1461
x"06c30",-- 1731
x"08340",-- 2100
x"09b00",-- 2480
x"0b670",-- 2919
x"0d0b0",-- 3339
x"0eb10",-- 3761
x"10840",-- 4228
x"12250",-- 4645
x"13bf0",-- 5055
x"14750",-- 5237
x"15220",-- 5410
x"15120",-- 5394
x"14af0",-- 5295
x"13580",-- 4952
x"10c30",-- 4291
x"0e040",-- 3588
x"0a640",-- 2660
x"06c70",-- 1735
x"01f90",-- 505
x"fd3b0",-- -709
x"f8610",-- -1951
x"f3f30",-- -3085
x"efed0",-- -4115
x"ebd80",-- -5160
x"e8b70",-- -5961
x"e63d0",-- -6595
x"e5200",-- -6880
x"e4940",-- -7020
x"e4d80",-- -6952
x"e61e0",-- -6626
x"e83f0",-- -6081
x"eb470",-- -5305
x"eeaf0",-- -4433
x"f29d0",-- -3427
x"f6a00",-- -2400
x"fae30",-- -1309
x"fee80",-- -280
x"02a00",-- 672
x"05f90",-- 1529
x"08a40",-- 2212
x"0ad60",-- 2774
x"0c180",-- 3096
x"0cfe0",-- 3326
x"0cfc0",-- 3324
x"0c7f0",-- 3199
x"0b300",-- 2864
x"099e0",-- 2462
x"07c70",-- 1991
x"05b50",-- 1461
x"03650",-- 869
x"00fa0",-- 250
x"feee0",-- -274
x"fce10",-- -799
x"fb420",-- -1214
x"f9740",-- -1676
x"f8530",-- -1965
x"f75c0",-- -2212
x"f6f70",-- -2313
x"f6bb0",-- -2373
x"f6980",-- -2408
x"f6fd0",-- -2307
x"f7660",-- -2202
x"f8480",-- -1976
x"f8f70",-- -1801
x"f9e70",-- -1561
x"fad20",-- -1326
x"fbf90",-- -1031
x"fd060",-- -762
x"fe0f0",-- -497
x"ff380",-- -200
x"00250",-- 37
x"01380",-- 312
x"022a0",-- 554
x"03400",-- 832
x"040d0",-- 1037
x"04f50",-- 1269
x"057c0",-- 1404
x"06140",-- 1556
x"068c0",-- 1676
x"06d60",-- 1750
x"06e30",-- 1763
x"06760",-- 1654
x"05e40",-- 1508
x"04f00",-- 1264
x"04350",-- 1077
x"02670",-- 615
x"00cf0",-- 207
x"fe930",-- -365
x"fcd00",-- -816
x"faf50",-- -1291
x"f8a20",-- -1886
x"f7160",-- -2282
x"f4e90",-- -2839
x"f4750",-- -2955
x"f3560",-- -3242
x"f30e0",-- -3314
x"f2f80",-- -3336
x"f34d0",-- -3251
x"f4c30",-- -2877
x"f5ae0",-- -2642
x"f7900",-- -2160
x"f9100",-- -1776
x"fb240",-- -1244
x"fd470",-- -697
x"ff260",-- -218
x"00de0",-- 222
x"02640",-- 612
x"03b00",-- 944
x"04c20",-- 1218
x"05630",-- 1379
x"05ec0",-- 1516
x"05f80",-- 1528
x"05d60",-- 1494
x"05ab0",-- 1451
x"05530",-- 1363
x"051d0",-- 1309
x"04b80",-- 1208
x"04550",-- 1109
x"04370",-- 1079
x"04520",-- 1106
x"04840",-- 1156
x"04af0",-- 1199
x"04f20",-- 1266
x"05ae0",-- 1454
x"06610",-- 1633
x"074a0",-- 1866
x"07e20",-- 2018
x"08c00",-- 2240
x"09ee0",-- 2542
x"0b4a0",-- 2890
x"0c860",-- 3206
x"0d970",-- 3479
x"0ef20",-- 3826
x"10550",-- 4181
x"118b0",-- 4491
x"122f0",-- 4655
x"12520",-- 4690
x"122f0",-- 4655
x"11e20",-- 4578
x"10a90",-- 4265
x"0ea20",-- 3746
x"0c080",-- 3080
x"095d0",-- 2397
x"06050",-- 1541
x"02620",-- 610
x"fe430",-- -445
x"fa2f0",-- -1489
x"f67b0",-- -2437
x"f2b90",-- -3399
x"ef470",-- -4281
x"ec100",-- -5104
x"e9ef0",-- -5649
x"e8260",-- -6106
x"e75e0",-- -6306
x"e7100",-- -6384
x"e7c50",-- -6203
x"e9330",-- -5837
x"eb420",-- -5310
x"ede80",-- -4632
x"f0de0",-- -3874
x"f4710",-- -2959
x"f7fe0",-- -2050
x"fba30",-- -1117
x"fee10",-- -287
x"024b0",-- 587
x"05100",-- 1296
x"07670",-- 1895
x"090b0",-- 2315
x"0a430",-- 2627
x"0af70",-- 2807
x"0aeb0",-- 2795
x"0a5e0",-- 2654
x"09350",-- 2357
x"08230",-- 2083
x"06840",-- 1668
x"04bb0",-- 1211
x"02b70",-- 695
x"00e40",-- 228
x"ff560",-- -170
x"fdda0",-- -550
x"fc800",-- -896
x"fb520",-- -1198
x"faa30",-- -1373
x"fa550",-- -1451
x"fa0d0",-- -1523
x"f9ea0",-- -1558
x"fa080",-- -1528
x"fa580",-- -1448
x"facf0",-- -1329
x"fb220",-- -1246
x"fb9e0",-- -1122
x"fbfe0",-- -1026
x"fc8a0",-- -886
x"fcfa0",-- -774
x"fd670",-- -665
x"fdce0",-- -562
x"fe620",-- -414
x"fec10",-- -319
x"ff380",-- -200
x"ffd50",-- -43
x"00750",-- 117
x"01180",-- 280
x"01b00",-- 432
x"026b0",-- 619
x"02e00",-- 736
x"03710",-- 881
x"03ae0",-- 942
x"03e00",-- 992
x"03f10",-- 1009
x"03a80",-- 936
x"02e00",-- 736
x"02690",-- 617
x"01540",-- 340
x"00910",-- 145
x"fed50",-- -299
x"fd8d0",-- -627
x"fc640",-- -924
x"faf30",-- -1293
x"fa440",-- -1468
x"f8570",-- -1961
x"f80c0",-- -2036
x"f73e0",-- -2242
x"f7290",-- -2263
x"f6e10",-- -2335
x"f6820",-- -2430
x"f7470",-- -2233
x"f7a20",-- -2142
x"f8a70",-- -1881
x"f92a0",-- -1750
x"fa1b0",-- -1509
x"fb330",-- -1229
x"fc850",-- -891
x"fd680",-- -664
x"fe890",-- -375
x"ff790",-- -135
x"00850",-- 133
x"01630",-- 355
x"023a0",-- 570
x"030e0",-- 782
x"037b0",-- 891
x"042b0",-- 1067
x"048e0",-- 1166
x"05290",-- 1321
x"05ab0",-- 1451
x"05f30",-- 1523
x"06320",-- 1586
x"06810",-- 1665
x"07060",-- 1798
x"075d0",-- 1885
x"078d0",-- 1933
x"07c70",-- 1991
x"08490",-- 2121
x"08c20",-- 2242
x"094c0",-- 2380
x"09a90",-- 2473
x"0a4f0",-- 2639
x"0b510",-- 2897
x"0c3e0",-- 3134
x"0d400",-- 3392
x"0dfb0",-- 3579
x"0f180",-- 3864
x"0fd00",-- 4048
x"103b0",-- 4155
x"106b0",-- 4203
x"102c0",-- 4140
x"0f9c0",-- 3996
x"0e820",-- 3714
x"0cdc0",-- 3292
x"0ac30",-- 2755
x"08770",-- 2167
x"05a90",-- 1449
x"02750",-- 629
x"fefd0",-- -259
x"fbbd0",-- -1091
x"f8640",-- -1948
x"f4fa0",-- -2822
x"f1d40",-- -3628
x"eefd0",-- -4355
x"ece40",-- -4892
x"eb1d0",-- -5347
x"e9fc0",-- -5636
x"e9450",-- -5819
x"e9650",-- -5787
x"ea4e0",-- -5554
x"eb920",-- -5230
x"ed4f0",-- -4785
x"ef980",-- -4200
x"f2570",-- -3497
x"f5450",-- -2747
x"f8520",-- -1966
x"fb310",-- -1231
x"fe250",-- -475
x"00c80",-- 200
x"034e0",-- 846
x"052b0",-- 1323
x"06b30",-- 1715
x"07d00",-- 2000
x"08680",-- 2152
x"08b60",-- 2230
x"08730",-- 2163
x"080c0",-- 2060
x"072b0",-- 1835
x"063f0",-- 1599
x"051d0",-- 1309
x"03ea0",-- 1002
x"02c60",-- 710
x"019c0",-- 412
x"007d0",-- 125
x"ff920",-- -110
x"fec60",-- -314
x"fe0f0",-- -497
x"fd790",-- -647
x"fcf30",-- -781
x"fccd0",-- -819
x"fc960",-- -874
x"fc9b0",-- -869
x"fc780",-- -904
x"fc800",-- -896
x"fcb40",-- -844
x"fcda0",-- -806
x"fd270",-- -729
x"fd440",-- -700
x"fd8b0",-- -629
x"fddf0",-- -545
x"fe320",-- -462
x"fe890",-- -375
x"feb20",-- -334
x"ff010",-- -255
x"ff270",-- -217
x"ff680",-- -152
x"ff950",-- -107
x"ffad0",-- -83
x"ffea0",-- -22
x"ffcc0",-- -52
x"00020",-- 2
x"00120",-- 18
x"003e0",-- 62
x"00120",-- 18
x"fffd0",-- -3
x"fffb0",-- -5
x"ffe40",-- -28
x"ffbc0",-- -68
x"ff3a0",-- -198
x"fee90",-- -279
x"fe940",-- -364
x"fe870",-- -377
x"fdf30",-- -525
x"fd620",-- -670
x"fcc00",-- -832
x"fc6e0",-- -914
x"fc210",-- -991
x"fba40",-- -1116
x"fb4a0",-- -1206
x"faf00",-- -1296
x"fb020",-- -1278
x"fb1d0",-- -1251
x"fb240",-- -1244
x"fb480",-- -1208
x"fbae0",-- -1106
x"fc200",-- -992
x"fca80",-- -856
x"fd2e0",-- -722
x"fdc40",-- -572
x"fe530",-- -429
x"ff110",-- -239
x"ffce0",-- -50
x"007b0",-- 123
x"013b0",-- 315
x"01e00",-- 480
x"02a70",-- 679
x"03790",-- 889
x"04620",-- 1122
x"051a0",-- 1306
x"05bc0",-- 1468
x"06810",-- 1665
x"075b0",-- 1883
x"08280",-- 2088
x"08d70",-- 2263
x"09790",-- 2425
x"0a110",-- 2577
x"0abe0",-- 2750
x"0b5b0",-- 2907
x"0bd60",-- 3030
x"0c340",-- 3124
x"0cf50",-- 3317
x"0d830",-- 3459
x"0e1e0",-- 3614
x"0e9b0",-- 3739
x"0ee00",-- 3808
x"0f360",-- 3894
x"0f1f0",-- 3871
x"0f400",-- 3904
x"0e980",-- 3736
x"0dd60",-- 3542
x"0cc80",-- 3272
x"0b400",-- 2880
x"09b70",-- 2487
x"07710",-- 1905
x"050e0",-- 1294
x"022b0",-- 555
x"ff8d0",-- -115
x"fca30",-- -861
x"f9940",-- -1644
x"f69b0",-- -2405
x"f3c20",-- -3134
x"f17f0",-- -3713
x"ef5e0",-- -4258
x"edba0",-- -4678
x"ec3f0",-- -5057
x"eba90",-- -5207
x"eb8e0",-- -5234
x"ec030",-- -5117
x"ecd50",-- -4907
x"edfb0",-- -4613
x"efc70",-- -4153
x"f1c00",-- -3648
x"f4200",-- -3040
x"f6620",-- -2462
x"f8cd0",-- -1843
x"fb250",-- -1243
x"fd790",-- -647
x"ff900",-- -112
x"01560",-- 342
x"02d90",-- 729
x"041c0",-- 1052
x"051a0",-- 1306
x"05d80",-- 1496
x"06440",-- 1604
x"06580",-- 1624
x"06500",-- 1616
x"06160",-- 1558
x"05c70",-- 1479
x"05440",-- 1348
x"04ae0",-- 1198
x"04030",-- 1027
x"036d0",-- 877
x"02dc0",-- 732
x"022f0",-- 559
x"01990",-- 409
x"01220",-- 290
x"00b20",-- 178
x"00570",-- 87
x"000c0",-- 12
x"ffb00",-- -80
x"ff6a0",-- -150
x"ff2e0",-- -210
x"ff1f0",-- -225
x"feee0",-- -274
x"febb0",-- -325
x"fe9b0",-- -357
x"fe7a0",-- -390
x"fe5d0",-- -419
x"fe3c0",-- -452
x"fe170",-- -489
x"fdfd0",-- -515
x"fdd10",-- -559
x"fdb70",-- -585
x"fdd00",-- -560
x"fd970",-- -617
x"fd940",-- -620
x"fd6d0",-- -659
x"fd5e0",-- -674
x"fd810",-- -639
x"fd880",-- -632
x"fd990",-- -615
x"fd8b0",-- -629
x"fd9c0",-- -612
x"fdb20",-- -590
x"fdae0",-- -594
x"fdab0",-- -597
x"fd940",-- -620
x"fd800",-- -640
x"fdb80",-- -584
x"fdce0",-- -562
x"fdd50",-- -555
x"fdd10",-- -559
x"fdce0",-- -562
x"fe210",-- -479
x"fe120",-- -494
x"fe3c0",-- -452
x"fe3f0",-- -449
x"fe5f0",-- -417
x"fe960",-- -362
x"fea80",-- -344
x"fea30",-- -349
x"fea70",-- -345
x"febc0",-- -324
x"fecb0",-- -309
x"feca0",-- -310
x"fec80",-- -312
x"fec80",-- -312
x"fecb0",-- -309
x"ff0c0",-- -244
x"ff2b0",-- -213
x"ff760",-- -138
x"ffd60",-- -42
x"00320",-- 50
x"00af0",-- 175
x"013d0",-- 317
x"01f90",-- 505
x"02a20",-- 674
x"034f0",-- 847
x"04300",-- 1072
x"04fe0",-- 1278
x"05d50",-- 1493
x"06930",-- 1683
x"07510",-- 1873
x"08250",-- 2085
x"08f40",-- 2292
x"09d50",-- 2517
x"0a730",-- 2675
x"0b4f0",-- 2895
x"0c220",-- 3106
x"0cf70",-- 3319
x"0dd00",-- 3536
x"0e7d0",-- 3709
x"0f080",-- 3848
x"0f650",-- 3941
x"0fbd0",-- 4029
x"0fa40",-- 4004
x"0f580",-- 3928
x"0e950",-- 3733
x"0d8d0",-- 3469
x"0c460",-- 3142
x"0aa70",-- 2727
x"08a20",-- 2210
x"063a0",-- 1594
x"03db0",-- 987
x"01420",-- 322
x"fea50",-- -347
x"fbc70",-- -1081
x"f9160",-- -1770
x"f6a50",-- -2395
x"f4690",-- -2967
x"f2840",-- -3452
x"f0c80",-- -3896
x"ef8e0",-- -4210
x"eec80",-- -4408
x"ee6c0",-- -4500
x"ee620",-- -4510
x"ee9b0",-- -4453
x"ef3e0",-- -4290
x"f0480",-- -4024
x"f17f0",-- -3713
x"f2ee0",-- -3346
x"f4700",-- -2960
x"f5f30",-- -2573
x"f7a80",-- -2136
x"f9480",-- -1720
x"fae60",-- -1306
x"fc580",-- -936
x"fdae0",-- -594
x"fef70",-- -265
x"000c0",-- 12
x"01080",-- 264
x"01bd0",-- 445
x"02690",-- 617
x"02e00",-- 736
x"03450",-- 837
x"03970",-- 919
x"03b80",-- 952
x"03c90",-- 969
x"03cc0",-- 972
x"03d50",-- 981
x"03d00",-- 976
x"03ba0",-- 954
x"03900",-- 912
x"037c0",-- 892
x"03560",-- 854
x"032c0",-- 812
x"03040",-- 772
x"02b90",-- 697
x"02850",-- 645
x"024b0",-- 587
x"02000",-- 512
x"01bd0",-- 445
x"01620",-- 354
x"011f0",-- 287
x"00dc0",-- 220
x"00780",-- 120
x"fffe0",-- -2
x"ff8a0",-- -118
x"ff130",-- -237
x"feaf0",-- -337
x"fe3c0",-- -452
x"fdc20",-- -574
x"fd710",-- -655
x"fcf30",-- -781
x"fca80",-- -856
x"fc440",-- -956
x"fbf30",-- -1037
x"fbcb0",-- -1077
x"fb880",-- -1144
x"fb880",-- -1144
x"fb5c0",-- -1188
x"fb650",-- -1179
x"fb8b0",-- -1141
x"fbc10",-- -1087
x"fc250",-- -987
x"fc6e0",-- -914
x"fcc60",-- -826
x"fd330",-- -717
x"fda60",-- -602
x"fe300",-- -464
x"fea80",-- -344
x"ff070",-- -249
x"ff620",-- -158
x"ff9f0",-- -97
x"ffdd0",-- -35
x"fffe0",-- -2
x"fff30",-- -13
x"ffd60",-- -42
x"ff900",-- -112
x"ff4a0",-- -182
x"fef50",-- -267
x"fe8c0",-- -372
x"fe390",-- -455
x"fdfd0",-- -515
x"fdee0",-- -530
x"fdd50",-- -555
x"fdce0",-- -562
x"fde90",-- -535
x"fe0d0",-- -499
x"fe660",-- -410
x"fec60",-- -314
x"ff330",-- -205
x"ffc70",-- -57
x"006e0",-- 110
x"01330",-- 307
x"02070",-- 519
x"02d20",-- 722
x"03a80",-- 936
x"04800",-- 1152
x"05600",-- 1376
x"062b0",-- 1579
x"06e00",-- 1760
x"07970",-- 1943
x"08550",-- 2133
x"090e0",-- 2318
x"09bd0",-- 2493
x"0a680",-- 2664
x"0b100",-- 2832
x"0bcb0",-- 3019
x"0c780",-- 3192
x"0d1c0",-- 3356
x"0d860",-- 3462
x"0deb0",-- 3563
x"0e360",-- 3638
x"0e480",-- 3656
x"0e270",-- 3623
x"0db30",-- 3507
x"0cff0",-- 3327
x"0c0c0",-- 3084
x"0aea0",-- 2794
x"09670",-- 2407
x"07b00",-- 1968
x"05d00",-- 1488
x"03c20",-- 962
x"018d0",-- 397
x"ff400",-- -192
x"fd090",-- -759
x"fae60",-- -1306
x"f9060",-- -1786
x"f7430",-- -2237
x"f5b80",-- -2632
x"f4710",-- -2959
x"f3750",-- -3211
x"f2ca0",-- -3382
x"f25f0",-- -3489
x"f2410",-- -3519
x"f2550",-- -3499
x"f2a50",-- -3419
x"f3240",-- -3292
x"f3cf0",-- -3121
x"f48e0",-- -2930
x"f5660",-- -2714
x"f6500",-- -2480
x"f74d0",-- -2227
x"f84b0",-- -1973
x"f9330",-- -1741
x"fa190",-- -1511
x"fae10",-- -1311
x"fbbd0",-- -1091
x"fc8e0",-- -882
x"fd3f0",-- -705
x"fde70",-- -537
x"fe820",-- -382
x"ff180",-- -232
x"ffad0",-- -83
x"002a0",-- 42
x"008f0",-- 143
x"00f90",-- 249
x"01630",-- 355
x"01c60",-- 454
x"02110",-- 529
x"024b0",-- 587
x"027b0",-- 635
x"02b60",-- 694
x"02e00",-- 736
x"02e80",-- 744
x"02f40",-- 756
x"02dc0",-- 732
x"02d90",-- 729
x"02be0",-- 702
x"02990",-- 665
x"02670",-- 615
x"02030",-- 515
x"01c20",-- 450
x"016d0",-- 365
x"01180",-- 280
x"00b40",-- 180
x"00480",-- 72
x"ffea0",-- -22
x"ff8a0",-- -118
x"ff5d0",-- -163
x"fefd0",-- -259
x"fe7f0",-- -385
x"fe4d0",-- -435
x"fe050",-- -507
x"fddd0",-- -547
x"fd8d0",-- -627
x"fd270",-- -729
x"fd160",-- -746
x"fd040",-- -764
x"fd130",-- -749
x"fcf20",-- -782
x"fceb0",-- -789
x"fd2a0",-- -726
x"fd4c0",-- -692
x"fd920",-- -622
x"fd830",-- -637
x"fd9c0",-- -612
x"fdc40",-- -572
x"fdc10",-- -575
x"fdcc0",-- -564
x"fd990",-- -615
x"fd8d0",-- -627
x"fd800",-- -640
x"fd6a0",-- -662
x"fd5e0",-- -674
x"fd440",-- -700
x"fd270",-- -729
x"fd1b0",-- -741
x"fd150",-- -747
x"fd160",-- -746
x"fd180",-- -744
x"fd1d0",-- -739
x"fd380",-- -712
x"fd620",-- -670
x"fdae0",-- -594
x"fdf60",-- -522
x"fe3a0",-- -454
x"fea80",-- -344
x"ff350",-- -203
x"ffcc0",-- -52
x"004d0",-- 77
x"00de0",-- 222
x"01720",-- 370
x"02230",-- 547
x"02d40",-- 724
x"035e0",-- 862
x"03df0",-- 991
x"045d0",-- 1117
x"04e80",-- 1256
x"05680",-- 1384
x"05db0",-- 1499
x"06520",-- 1618
x"06c80",-- 1736
x"07630",-- 1891
x"07ec0",-- 2028
x"08820",-- 2178
x"09170",-- 2327
x"09bd0",-- 2493
x"0a7a0",-- 2682
x"0b240",-- 2852
x"0bba0",-- 3002
x"0c2d0",-- 3117
x"0c9a0",-- 3226
x"0cdc0",-- 3292
x"0ceb0",-- 3307
x"0cb80",-- 3256
x"0c480",-- 3144
x"0ba80",-- 2984
x"0ad60",-- 2774
x"09bc0",-- 2492
x"086e0",-- 2158
x"06ea0",-- 1770
x"05470",-- 1351
x"039c0",-- 924
x"01d50",-- 469
x"000a0",-- 10
x"fe4b0",-- -437
x"fcbe0",-- -834
x"fb4f0",-- -1201
x"f9fd0",-- -1539
x"f8d50",-- -1835
x"f7dd0",-- -2083
x"f7200",-- -2272
x"f6890",-- -2423
x"f6250",-- -2523
x"f5dd0",-- -2595
x"f5ba0",-- -2630
x"f5b30",-- -2637
x"f5d50",-- -2603
x"f6120",-- -2542
x"f65d0",-- -2467
x"f6bb0",-- -2373
x"f7290",-- -2263
x"f7a10",-- -2143
x"f82f0",-- -2001
x"f8c80",-- -1848
x"f95e0",-- -1698
x"f9fb0",-- -1541
x"faa70",-- -1369
x"fb570",-- -1193
x"fbf10",-- -1039
x"fc710",-- -911
x"fce40",-- -796
x"fd580",-- -680
x"fdb30",-- -589
x"fe0a0",-- -502
x"fe520",-- -430
x"fe9e0",-- -354
x"fef00",-- -272
x"ff3a0",-- -198
x"ff860",-- -122
x"ffce0",-- -50
x"00070",-- 7
x"00320",-- 50
x"006c0",-- 108
x"00990",-- 153
x"00c10",-- 193
x"00e60",-- 230
x"00f90",-- 249
x"01100",-- 272
x"011d0",-- 285
x"01270",-- 295
x"01350",-- 309
x"013b0",-- 315
x"01400",-- 320
x"01470",-- 327
x"01470",-- 327
x"013b0",-- 315
x"01180",-- 280
x"00fe0",-- 254
x"00f50",-- 245
x"00c50",-- 197
x"00870",-- 135
x"00520",-- 82
x"002b0",-- 43
x"00030",-- 3
x"ffe20",-- -30
x"ffad0",-- -83
x"ff8a0",-- -118
x"ff720",-- -142
x"ff490",-- -183
x"ff1f0",-- -225
x"fef00",-- -272
x"feca0",-- -310
x"fe910",-- -367
x"fe500",-- -432
x"fe140",-- -492
x"fdd30",-- -557
x"fda10",-- -607
x"fd710",-- -655
x"fd470",-- -697
x"fd1b0",-- -741
x"fd020",-- -766
x"fce90",-- -791
x"fccd0",-- -819
x"fccb0",-- -821
x"fcd00",-- -816
x"fcda0",-- -806
x"fce10",-- -799
x"fcf30",-- -781
x"fd150",-- -747
x"fd3b0",-- -709
x"fd6f0",-- -657
x"fd9c0",-- -612
x"fdd50",-- -555
x"fe200",-- -480
x"fe730",-- -397
x"feca0",-- -310
x"ff1f0",-- -225
x"ff8d0",-- -115
x"00000",-- 0
x"00640",-- 100
x"00d50",-- 213
x"013a0",-- 314
x"01ad0",-- 429
x"02260",-- 550
x"029e0",-- 670
x"031d0",-- 797
x"038a0",-- 906
x"04170",-- 1047
x"04a00",-- 1184
x"052b0",-- 1323
x"05c40",-- 1476
x"06430",-- 1603
x"06dc0",-- 1756
x"07740",-- 1908
x"081e0",-- 2078
x"08c20",-- 2242
x"095e0",-- 2398
x"0a140",-- 2580
x"0aa00",-- 2720
x"0b300",-- 2864
x"0b940",-- 2964
x"0be20",-- 3042
x"0c130",-- 3091
x"0c080",-- 3080
x"0bd00",-- 3024
x"0b6a0",-- 2922
x"0ad70",-- 2775
x"0a0d0",-- 2573
x"09130",-- 2323
x"07e40",-- 2020
x"06a50",-- 1701
x"05420",-- 1346
x"03da0",-- 986
x"02520",-- 594
x"00dc0",-- 220
x"ff800",-- -128
x"fe2a0",-- -470
x"fcf70",-- -777
x"fbd60",-- -1066
x"fadf0",-- -1313
x"fa110",-- -1519
x"f9660",-- -1690
x"f8d20",-- -1838
x"f8570",-- -1961
x"f80a0",-- -2038
x"f7d60",-- -2090
x"f7bf0",-- -2113
x"f7c90",-- -2103
x"f7e00",-- -2080
x"f8190",-- -2023
x"f8780",-- -1928
x"f8da0",-- -1830
x"f94a0",-- -1718
x"f9bc0",-- -1604
x"fa2a0",-- -1494
x"fa820",-- -1406
x"fac50",-- -1339
x"fade0",-- -1314
x"fadf0",-- -1313
x"fae60",-- -1306
x"faed0",-- -1299
x"fb0e0",-- -1266
x"fb450",-- -1211
x"fb880",-- -1144
x"fbd00",-- -1072
x"fc340",-- -972
x"fc930",-- -877
x"fce90",-- -791
x"fd380",-- -712
x"fd830",-- -637
x"fdb30",-- -589
x"fde70",-- -537
x"fe320",-- -462
x"fe750",-- -395
x"fec60",-- -314
x"ff0b0",-- -245
x"ff600",-- -160
x"ffb80",-- -72
x"fff90",-- -7
x"003e0",-- 62
x"00870",-- 135
x"00c00",-- 192
x"00f20",-- 242
x"01180",-- 280
x"01310",-- 305
x"01420",-- 322
x"01440",-- 324
x"014f0",-- 335
x"01650",-- 357
x"015e0",-- 350
x"01580",-- 344
x"015d0",-- 349
x"01650",-- 357
x"015d0",-- 349
x"01470",-- 327
x"01310",-- 305
x"010e0",-- 270
x"00e90",-- 233
x"00c10",-- 193
x"00820",-- 130
x"00410",-- 65
x"fffb0",-- -5
x"ffb80",-- -72
x"ff710",-- -143
x"ff240",-- -220
x"fede0",-- -290
x"fea50",-- -347
x"fe750",-- -395
x"fe3e0",-- -450
x"fe210",-- -479
x"fdf10",-- -527
x"fdd60",-- -554
x"fdbc0",-- -580
x"fdb30",-- -589
x"fda30",-- -605
x"fd8b0",-- -629
x"fd880",-- -632
x"fd860",-- -634
x"fd950",-- -619
x"fda80",-- -600
x"fdb00",-- -592
x"fdc40",-- -572
x"fdf10",-- -527
x"fe1b0",-- -485
x"fe490",-- -439
x"fe820",-- -382
x"fec10",-- -319
x"ff060",-- -250
x"ff540",-- -172
x"ff9f0",-- -97
x"fff10",-- -15
x"003e0",-- 62
x"00990",-- 153
x"01010",-- 257
x"017b0",-- 379
x"01f60",-- 502
x"02750",-- 629
x"02fe0",-- 766
x"037b0",-- 891
x"04140",-- 1044
x"04ac0",-- 1196
x"05470",-- 1351
x"05e50",-- 1509
x"068b0",-- 1675
x"073a0",-- 1850
x"07ef0",-- 2031
x"089a0",-- 2202
x"094c0",-- 2380
x"09ee0",-- 2542
x"0a750",-- 2677
x"0aef0",-- 2799
x"0b350",-- 2869
x"0b650",-- 2917
x"0b5e0",-- 2910
x"0b310",-- 2865
x"0ae10",-- 2785
x"0a4f0",-- 2639
x"09940",-- 2452
x"08a00",-- 2208
x"079c0",-- 1948
x"067a0",-- 1658
x"05400",-- 1344
x"03ea0",-- 1002
x"027f0",-- 639
x"012c0",-- 300
x"ffe90",-- -23
x"feb60",-- -330
x"fd810",-- -639
x"fc760",-- -906
x"fb920",-- -1134
x"facf0",-- -1329
x"fa370",-- -1481
x"f9ad0",-- -1619
x"f9480",-- -1720
x"f9150",-- -1771
x"f8f20",-- -1806
x"f9040",-- -1788
x"f9240",-- -1756
x"f9660",-- -1690
x"f9bc0",-- -1604
x"fa050",-- -1531
x"fa6b0",-- -1429
x"faad0",-- -1363
x"faca0",-- -1334
x"fad40",-- -1324
x"fab90",-- -1351
x"fa9b0",-- -1381
x"fa710",-- -1423
x"fa550",-- -1451
x"fa4b0",-- -1461
x"fa520",-- -1454
x"fa7d0",-- -1411
x"faaf0",-- -1361
x"faee0",-- -1298
x"fb150",-- -1259
x"fb470",-- -1209
x"fb740",-- -1164
x"fba30",-- -1117
x"fbd00",-- -1072
x"fbfe0",-- -1026
x"fc340",-- -972
x"fc820",-- -894
x"fce80",-- -792
x"fd380",-- -712
x"fd9f0",-- -609
x"fe070",-- -505
x"fe7f0",-- -385
x"fee10",-- -287
x"ff3b0",-- -197
x"ff860",-- -122
x"ffb70",-- -73
x"fff30",-- -13
x"00230",-- 35
x"00430",-- 67
x"005d0",-- 93
x"00800",-- 128
x"00a80",-- 168
x"00cf0",-- 207
x"00f40",-- 244
x"01170",-- 279
x"013d0",-- 317
x"01600",-- 352
x"016a0",-- 362
x"017c0",-- 380
x"017b0",-- 379
x"015e0",-- 350
x"014a0",-- 330
x"011a0",-- 282
x"00e10",-- 225
x"00a80",-- 168
x"00620",-- 98
x"00250",-- 37
x"fff80",-- -8
x"ffb20",-- -78
x"ff760",-- -138
x"ff4f0",-- -177
x"ff1d0",-- -227
x"fefa0",-- -262
x"fee10",-- -287
x"fec80",-- -312
x"fead0",-- -339
x"fe8f0",-- -369
x"fe820",-- -382
x"fe7b0",-- -389
x"fe660",-- -410
x"fe5a0",-- -422
x"fe570",-- -425
x"fe4d0",-- -435
x"fe460",-- -442
x"fe480",-- -440
x"fe490",-- -439
x"fe4b0",-- -437
x"fe5f0",-- -417
x"fe620",-- -414
x"fe820",-- -382
x"feb40",-- -332
x"fed40",-- -300
x"ff060",-- -250
x"ff510",-- -175
x"ff940",-- -108
x"ffe40",-- -28
x"003a0",-- 58
x"009e0",-- 158
x"01150",-- 277
x"01970",-- 407
x"020c0",-- 524
x"02890",-- 649
x"03130",-- 787
x"039c0",-- 924
x"04260",-- 1062
x"04b60",-- 1206
x"054a0",-- 1354
x"05e50",-- 1509
x"06840",-- 1668
x"071c0",-- 1820
x"07c60",-- 1990
x"08640",-- 2148
x"09080",-- 2312
x"09a30",-- 2467
x"0a200",-- 2592
x"0a810",-- 2689
x"0ac50",-- 2757
x"0ad40",-- 2772
x"0ab10",-- 2737
x"0a630",-- 2659
x"09db0",-- 2523
x"09290",-- 2345
x"08440",-- 2116
x"07450",-- 1861
x"060f0",-- 1551
x"04d10",-- 1233
x"03830",-- 899
x"02110",-- 529
x"00a80",-- 168
x"ff4f0",-- -177
x"fe0a0",-- -502
x"fced0",-- -787
x"fbe00",-- -1056
x"faf20",-- -1294
x"fa480",-- -1464
x"f9c60",-- -1594
x"f9740",-- -1676
x"f9420",-- -1726
x"f9360",-- -1738
x"f9660",-- -1690
x"f9a30",-- -1629
x"f9f10",-- -1551
x"fa500",-- -1456
x"fab20",-- -1358
x"fb130",-- -1261
x"fb650",-- -1179
x"fb860",-- -1146
x"fb760",-- -1162
x"fb520",-- -1198
x"fb2c0",-- -1236
x"fb070",-- -1273
x"fae30",-- -1309
x"fadc0",-- -1316
x"fadf0",-- -1313
x"faf20",-- -1294
x"fb0e0",-- -1266
x"fb240",-- -1244
x"fb480",-- -1208
x"fb620",-- -1182
x"fb680",-- -1176
x"fb8d0",-- -1139
x"fbae0",-- -1106
x"fbd00",-- -1072
x"fc070",-- -1017
x"fc350",-- -971
x"fc7b0",-- -901
x"fccd0",-- -819
x"fd1d0",-- -739
x"fd7b0",-- -645
x"fdd80",-- -552
x"fe320",-- -462
x"fe8a0",-- -374
x"fed90",-- -295
x"ff070",-- -249
x"ff310",-- -207
x"ff5b0",-- -165
x"ff950",-- -107
x"ffc90",-- -55
x"fff30",-- -13
x"00210",-- 33
x"004e0",-- 78
x"00870",-- 135
x"00c60",-- 198
x"00ed0",-- 237
x"01150",-- 277
x"013f0",-- 319
x"01440",-- 324
x"01380",-- 312
x"01180",-- 280
x"00fe0",-- 254
x"00cb0",-- 203
x"009d0",-- 157
x"00660",-- 102
x"00350",-- 53
x"00030",-- 3
x"ffcb0",-- -53
x"ffae0",-- -82
x"ff850",-- -123
x"ff740",-- -140
x"ff580",-- -168
x"ff3d0",-- -195
x"ff310",-- -207
x"ff240",-- -220
x"ff1a0",-- -230
x"ff0e0",-- -242
x"ff070",-- -249
x"fef30",-- -269
x"fee40",-- -284
x"fede0",-- -290
x"fed70",-- -297
x"febb0",-- -325
x"feaf0",-- -337
x"fea20",-- -350
x"fea80",-- -344
x"feaa0",-- -342
x"feaf0",-- -337
x"fed40",-- -300
x"fef00",-- -272
x"ff1f0",-- -225
x"ff470",-- -185
x"ff710",-- -143
x"ffbc0",-- -68
x"fffb0",-- -5
x"00480",-- 72
x"00a70",-- 167
x"01080",-- 264
x"01810",-- 385
x"01ef0",-- 495
x"02780",-- 632
x"03090",-- 777
x"03a80",-- 936
x"043c0",-- 1084
x"04d90",-- 1241
x"05900",-- 1424
x"063e0",-- 1598
x"07080",-- 1800
x"07d00",-- 2000
x"08b30",-- 2227
x"09920",-- 2450
x"0a640",-- 2660
x"0b060",-- 2822
x"0b8b0",-- 2955
x"0c080",-- 3080
x"0c430",-- 3139
x"0c3b0",-- 3131
x"0bcc0",-- 3020
x"0b2c0",-- 2860
x"0a680",-- 2664
x"09600",-- 2400
x"08120",-- 2066
x"06810",-- 1665
x"04e30",-- 1251
x"032e0",-- 814
x"01770",-- 375
x"ffa30",-- -93
x"fdd00",-- -560
x"fc2a0",-- -982
x"fac00",-- -1344
x"f9900",-- -1648
x"f87a0",-- -1926
x"f7a90",-- -2135
x"f7130",-- -2285
x"f6cf0",-- -2353
x"f6c10",-- -2367
x"f6eb0",-- -2325
x"f7330",-- -2253
x"f7b00",-- -2128
x"f8530",-- -1965
x"f90b0",-- -1781
x"f9d50",-- -1579
x"fa910",-- -1391
x"fb420",-- -1214
x"fbda0",-- -1062
x"fc5f0",-- -929
x"fcbc0",-- -836
x"fcff0",-- -769
x"fd100",-- -752
x"fd070",-- -761
x"fd0b0",-- -757
x"fd060",-- -762
x"fd090",-- -759
x"fcff0",-- -769
x"fcff0",-- -769
x"fd060",-- -762
x"fd130",-- -749
x"fd130",-- -749
x"fd020",-- -766
x"fce10",-- -799
x"fcbb0",-- -837
x"fcaa0",-- -854
x"fc9b0",-- -869
x"fc8a0",-- -886
x"fc780",-- -904
x"fc890",-- -887
x"fc990",-- -871
x"fcc80",-- -824
x"fcf20",-- -782
x"fd200",-- -736
x"fd6f0",-- -657
x"fdb50",-- -587
x"fe0f0",-- -497
x"fe690",-- -407
x"fecb0",-- -309
x"ff300",-- -208
x"ff950",-- -107
x"fff80",-- -8
x"005d0",-- 93
x"00c00",-- 192
x"010d0",-- 269
x"01360",-- 310
x"015b0",-- 347
x"017b0",-- 379
x"01770",-- 375
x"015e0",-- 350
x"012b0",-- 299
x"00f90",-- 249
x"00c80",-- 200
x"00930",-- 147
x"00460",-- 70
x"fff10",-- -15
x"ffd50",-- -43
x"ffb00",-- -80
x"ff8d0",-- -115
x"ff630",-- -157
x"ff440",-- -188
x"ff380",-- -200
x"ff2b0",-- -213
x"ff2b0",-- -213
x"ff150",-- -235
x"ff070",-- -249
x"ff020",-- -254
x"ff060",-- -250
x"fefd0",-- -259
x"fef00",-- -272
x"fef30",-- -269
x"ff070",-- -249
x"ff110",-- -239
x"ff180",-- -232
x"ff260",-- -218
x"ff350",-- -203
x"ff510",-- -175
x"ff6f0",-- -145
x"ffa30",-- -93
x"ffd50",-- -43
x"00140",-- 20
x"00690",-- 105
x"00cf0",-- 207
x"013b0",-- 315
x"01c20",-- 450
x"024e0",-- 590
x"02e30",-- 739
x"03810",-- 897
x"04370",-- 1079
x"05060",-- 1286
x"05c90",-- 1481
x"06930",-- 1683
x"076f0",-- 1903
x"08720",-- 2162
x"09770",-- 2423
x"0a8c0",-- 2700
x"0b9e0",-- 2974
x"0cbd0",-- 3261
x"0dec0",-- 3564
x"0ef70",-- 3831
x"0fbd0",-- 4029
x"100e0",-- 4110
x"10450",-- 4165
x"10160",-- 4118
x"0f6c0",-- 3948
x"0e480",-- 3656
x"0c950",-- 3221
x"0ab40",-- 2740
x"08810",-- 2177
x"06140",-- 1556
x"034f0",-- 847
x"00800",-- 128
x"fdd00",-- -560
x"fb390",-- -1223
x"f8eb0",-- -1813
x"f6940",-- -2412
x"f4a80",-- -2904
x"f3130",-- -3309
x"f1fb0",-- -3589
x"f1380",-- -3784
x"f0c00",-- -3904
x"f0ad0",-- -3923
x"f0e40",-- -3868
x"f1680",-- -3736
x"f2100",-- -3568
x"f3070",-- -3321
x"f3f60",-- -3082
x"f51b0",-- -2789
x"f6490",-- -2487
x"f78d0",-- -2163
x"f8f80",-- -1800
x"fa4d0",-- -1459
x"fbad0",-- -1107
x"fceb0",-- -789
x"fe570",-- -425
x"ffad0",-- -83
x"00f40",-- 244
x"02030",-- 515
x"02f70",-- 759
x"03d60",-- 982
x"046c0",-- 1132
x"04be0",-- 1214
x"04be0",-- 1214
x"048c0",-- 1164
x"04340",-- 1076
x"03950",-- 917
x"02b70",-- 695
x"01810",-- 385
x"004d0",-- 77
x"ff1a0",-- -230
x"fdd50",-- -555
x"fc730",-- -909
x"fb1a0",-- -1254
x"f9f10",-- -1551
x"f8fa0",-- -1798
x"f82b0",-- -2005
x"f78d0",-- -2163
x"f7330",-- -2253
x"f7450",-- -2235
x"f78e0",-- -2162
x"f81c0",-- -2020
x"f8f70",-- -1801
x"f9c90",-- -1591
x"faf20",-- -1294
x"fc0f0",-- -1009
x"fd4e0",-- -690
x"feac0",-- -340
x"ffdd0",-- -35
x"010e0",-- 270
x"01f30",-- 499
x"02f70",-- 759
x"03c10",-- 961
x"04570",-- 1111
x"04a70",-- 1191
x"04ae0",-- 1198
x"04cd0",-- 1229
x"04a90",-- 1193
x"045f0",-- 1119
x"03d60",-- 982
x"033a0",-- 826
x"029b0",-- 667
x"01d80",-- 472
x"01040",-- 260
x"00160",-- 22
x"ff180",-- -232
x"fe3a0",-- -454
x"fd6d0",-- -659
x"fcbb0",-- -837
x"fc070",-- -1017
x"fb6c0",-- -1172
x"fb330",-- -1229
x"fb240",-- -1244
x"fb520",-- -1198
x"fba40",-- -1116
x"fc1c0",-- -996
x"fcda0",-- -806
x"fdb50",-- -587
x"fecf0",-- -305
x"ffc90",-- -55
x"00c10",-- 193
x"01bd0",-- 445
x"02cc0",-- 716
x"03e50",-- 997
x"04db0",-- 1243
x"05b50",-- 1461
x"06640",-- 1636
x"07580",-- 1880
x"084d0",-- 2125
x"09450",-- 2373
x"0a4f0",-- 2639
x"0b3d0",-- 2877
x"0c5c0",-- 3164
x"0dad0",-- 3501
x"0f1c0",-- 3868
x"108e0",-- 4238
x"11d80",-- 4568
x"13150",-- 4885
x"145e0",-- 5214
x"15c40",-- 5572
x"16c70",-- 5831
x"17240",-- 5924
x"16b80",-- 5816
x"16050",-- 5637
x"149b0",-- 5275
x"129a0",-- 4762
x"0f590",-- 3929
x"0b810",-- 2945
x"07590",-- 1881
x"03180",-- 792
x"febb0",-- -325
x"f9f60",-- -1546
x"f5720",-- -2702
x"f14c0",-- -3764
x"ee0b0",-- -4597
x"eb360",-- -5322
x"e8df0",-- -5921
x"e72e0",-- -6354
x"e6420",-- -6590
x"e6490",-- -6583
x"e6aa0",-- -6486
x"e7d30",-- -6189
x"e92f0",-- -5841
x"eb040",-- -5372
x"ed180",-- -4840
x"ef7f0",-- -4225
x"f2010",-- -3583
x"f4960",-- -2922
x"f7270",-- -2265
x"f9a30",-- -1629
x"fc2d0",-- -979
x"febe0",-- -322
x"016d0",-- 365
x"038f0",-- 911
x"05a40",-- 1444
x"07770",-- 1911
x"09510",-- 2385
x"0ade0",-- 2782
x"0bc40",-- 3012
x"0c360",-- 3126
x"0c110",-- 3089
x"0bf30",-- 3059
x"0b330",-- 2867
x"09d80",-- 2520
x"07c20",-- 1986
x"05450",-- 1349
x"02c00",-- 704
x"00250",-- 37
x"fd800",-- -640
x"fa500",-- -1456
x"f7980",-- -2152
x"f5420",-- -2750
x"f3970",-- -3177
x"f2340",-- -3532
x"f1090",-- -3831
x"f0440",-- -4028
x"f0120",-- -4078
x"f0c60",-- -3898
x"f1790",-- -3719
x"f2b90",-- -3399
x"f3a60",-- -3162
x"f5290",-- -2775
x"f6e80",-- -2328
x"f8d70",-- -1833
x"facf0",-- -1329
x"fc050",-- -1019
x"fde70",-- -537
x"ff7c0",-- -132
x"01c60",-- 454
x"033d0",-- 829
x"04b90",-- 1209
x"05f10",-- 1521
x"07490",-- 1865
x"089d0",-- 2205
x"093d0",-- 2365
x"09b80",-- 2488
x"095d0",-- 2397
x"09330",-- 2355
x"08950",-- 2197
x"07990",-- 1945
x"05fb0",-- 1531
x"04390",-- 1081
x"025c0",-- 604
x"005a0",-- 90
x"fe890",-- -375
x"fcbe0",-- -834
x"fb1f0",-- -1249
x"f9480",-- -1720
x"f8500",-- -1968
x"f76b0",-- -2197
x"f7400",-- -2240
x"f7040",-- -2300
x"f6fa0",-- -2310
x"f7790",-- -2183
x"f8570",-- -1961
x"fa170",-- -1513
x"fb650",-- -1179
x"fd240",-- -732
x"ff090",-- -247
x"019f0",-- 415
x"04730",-- 1139
x"07350",-- 1845
x"09f80",-- 2552
x"0c540",-- 3156
x"0f2c0",-- 3884
x"11c10",-- 4545
x"146e0",-- 5230
x"16720",-- 5746
x"18a00",-- 6304
x"1a750",-- 6773
x"1cb40",-- 7348
x"1ed60",-- 7894
x"207a0",-- 8314
x"21ad0",-- 8621
x"22430",-- 8771
x"22e30",-- 8931
x"22050",-- 8709
x"205a0",-- 8282
x"1cb80",-- 7352
x"18110",-- 6161
x"120a0",-- 4618
x"0b770",-- 2935
x"03d50",-- 981
x"fb5e0",-- -1186
x"f35e0",-- -3234
x"ebb80",-- -5192
x"e54d0",-- -6835
x"df680",-- -8344
x"db1b0",-- -9445
x"d7e30",-- -10269
x"d65b0",-- -10661
x"d62b0",-- -10709
x"d72c0",-- -10452
x"d9340",-- -9932
x"dc060",-- -9210
x"dfce0",-- -8242
x"e3d40",-- -7212
x"e8940",-- -5996
x"ed6d0",-- -4755
x"f2d20",-- -3374
x"f7da0",-- -2086
x"fd100",-- -752
x"02230",-- 547
x"074a0",-- 1866
x"0c230",-- 3107
x"102d0",-- 4141
x"13dc0",-- 5084
x"16a90",-- 5801
x"19010",-- 6401
x"19ff0",-- 6655
x"1a0e0",-- 6670
x"18ac0",-- 6316
x"16700",-- 5744
x"13420",-- 4930
x"0f2b0",-- 3883
x"0a430",-- 2627
x"04a20",-- 1186
x"feee0",-- -274
x"f92c0",-- -1748
x"f3b60",-- -3146
x"ee6c0",-- -4500
x"e9cf0",-- -5681
x"e5ca0",-- -6710
x"e2f00",-- -7440
x"e1250",-- -7899
x"e03a0",-- -8134
x"e02b0",-- -8149
x"e1050",-- -7931
x"e34c0",-- -7348
x"e62b0",-- -6613
x"e9cc0",-- -5684
x"edc40",-- -4668
x"f2820",-- -3454
x"f7680",-- -2200
x"fcc60",-- -826
x"02080",-- 520
x"06a50",-- 1701
x"0b3f0",-- 2879
x"0f060",-- 3846
x"130e0",-- 4878
x"156f0",-- 5487
x"17550",-- 5973
x"17b40",-- 6068
x"17970",-- 6039
x"16c30",-- 5827
x"14dc0",-- 5340
x"121b0",-- 4635
x"0dfb0",-- 3579
x"0a120",-- 2578
x"058a0",-- 1418
x"01580",-- 344
x"fc760",-- -906
x"f80d0",-- -2035
x"f3f10",-- -3087
x"f0960",-- -3946
x"ee2d0",-- -4563
x"ec100",-- -5104
x"eaed0",-- -5395
x"e9f10",-- -5647
x"ea740",-- -5516
x"eb4a0",-- -5302
x"ed540",-- -4780
x"ef6a0",-- -4246
x"f24e0",-- -3506
x"f5470",-- -2745
x"f90e0",-- -1778
x"fd440",-- -700
x"014f0",-- 335
x"059e0",-- 1438
x"094e0",-- 2382
x"0d950",-- 3477
x"11180",-- 4376
x"14770",-- 5239
x"16c20",-- 5826
x"18700",-- 6256
x"199b0",-- 6555
x"19f10",-- 6641
x"19cd0",-- 6605
x"18900",-- 6288
x"17330",-- 5939
x"15a60",-- 5542
x"143e0",-- 5182
x"133a0",-- 4922
x"12b60",-- 4790
x"13120",-- 4882
x"14570",-- 5207
x"161d0",-- 5661
x"17e20",-- 6114
x"18be0",-- 6334
x"1a180",-- 6680
x"1ad60",-- 6870
x"19a30",-- 6563
x"155b0",-- 5467
x"0f530",-- 3923
x"08f00",-- 2288
x"01d60",-- 470
x"f9c70",-- -1593
x"f0490",-- -4023
x"e8260",-- -6106
x"e24e0",-- -7602
x"df0e0",-- -8434
x"dc7e0",-- -9090
x"daf30",-- -9485
x"db4f0",-- -9393
x"dd9d0",-- -8803
x"e1190",-- -7911
x"e42d0",-- -7123
x"e7150",-- -6379
x"ea2d0",-- -5587
x"edc90",-- -4663
x"f0de0",-- -3874
x"f4440",-- -3004
x"f8110",-- -2031
x"fc960",-- -874
x"01170",-- 279
x"061b0",-- 1563
x"0b830",-- 2947
x"10ef0",-- 4335
x"16370",-- 5687
x"198a0",-- 6538
x"1b0f0",-- 6927
x"1b210",-- 6945
x"1a340",-- 6708
x"16690",-- 5737
x"10590",-- 4185
x"08bd0",-- 2237
x"00ad0",-- 173
x"f8ff0",-- -1793
x"f1b80",-- -3656
x"eb240",-- -5340
x"e5ba0",-- -6726
x"e2b00",-- -7504
x"e1930",-- -7789
x"e1e70",-- -7705
x"e3250",-- -7387
x"e53b0",-- -6853
x"e71a0",-- -6374
x"e8aa0",-- -5974
x"ea7b0",-- -5509
x"ec6f0",-- -5009
x"ee990",-- -4455
x"f03e0",-- -4034
x"f28a0",-- -3446
x"f6520",-- -2478
x"fbdf0",-- -1057
x"026b0",-- 619
x"09580",-- 2392
x"0f9e0",-- 3998
x"15f00",-- 5616
x"1c000",-- 7168
x"20970",-- 8343
x"225c0",-- 8796
x"211f0",-- 8479
x"1db40",-- 7604
x"17500",-- 5968
x"10e60",-- 4326
x"09030",-- 2307
x"01540",-- 340
x"f9330",-- -1741
x"f31b0",-- -3301
x"efa10",-- -4191
x"ee3a0",-- -4550
x"ee0f0",-- -4593
x"ee240",-- -4572
x"ef390",-- -4295
x"f0820",-- -3966
x"f1ef0",-- -3601
x"f2620",-- -3486
x"f19c0",-- -3684
x"ef900",-- -4208
x"ef480",-- -4280
x"efdd0",-- -4131
x"f12e0",-- -3794
x"f3f80",-- -3080
x"f7f80",-- -2056
x"fdad0",-- -595
x"03dd0",-- 989
x"0af90",-- 2809
x"10a20",-- 4258
x"148c0",-- 5260
x"167f0",-- 5759
x"16cd0",-- 5837
x"14ed0",-- 5357
x"12500",-- 4688
x"0e950",-- 3733
x"0a190",-- 2585
x"065f0",-- 1631
x"042d0",-- 1069
x"040c0",-- 1036
x"04580",-- 1112
x"050e0",-- 1294
x"063a0",-- 1594
x"083f0",-- 2111
x"0abb0",-- 2747
x"0cf50",-- 3317
x"0e270",-- 3623
x"0f950",-- 3989
x"11a60",-- 4518
x"149a0",-- 5274
x"176c0",-- 5996
x"1ad90",-- 6873
x"1f320",-- 7986
x"22920",-- 8850
x"24d10",-- 9425
x"24ef0",-- 9455
x"23690",-- 9065
x"1f0a0",-- 7946
x"17330",-- 5939
x"0ba40",-- 2980
x"fefa0",-- -262
x"f31d0",-- -3299
x"e8690",-- -6039
x"ded20",-- -8494
x"d7020",-- -10494
x"d32a0",-- -11478
x"d2d50",-- -11563
x"d5590",-- -10919
x"d86c0",-- -10132
x"dbfc0",-- -9220
x"dfea0",-- -8214
x"e3e30",-- -7197
x"e7900",-- -6256
x"eada0",-- -5414
x"eeac0",-- -4436
x"f38e0",-- -3186
x"f9540",-- -1708
x"00490",-- 73
x"094c0",-- 2380
x"13010",-- 4865
x"1c390",-- 7225
x"23470",-- 9031
x"27ce0",-- 10190
x"296a0",-- 10602
x"27c10",-- 10177
x"21be0",-- 8638
x"17990",-- 6041
x"0b5d0",-- 2909
x"ff180",-- -232
x"f3840",-- -3196
x"e9480",-- -5816
x"e1840",-- -7804
x"dcd20",-- -9006
x"db8b0",-- -9333
x"dc9c0",-- -9060
x"df2c0",-- -8404
x"e20f0",-- -7665
x"e4b20",-- -6990
x"e6a00",-- -6496
x"e7480",-- -6328
x"e7d30",-- -6189
x"e8ab0",-- -5973
x"ea560",-- -5546
x"eca20",-- -4958
x"f1100",-- -3824
x"f8c30",-- -1853
x"02d20",-- 722
x"0d920",-- 3474
x"16c80",-- 5832
x"1f1e0",-- 7966
x"24c50",-- 9413
x"27c90",-- 10185
x"27530",-- 10067
x"22ab0",-- 8875
x"1b740",-- 7028
x"122c0",-- 4652
x"0a6d0",-- 2669
x"02780",-- 632
x"fb0e0",-- -1266
x"f6280",-- -2520
x"f34a0",-- -3254
x"f2050",-- -3579
x"f08f0",-- -3953
x"f0320",-- -4046
x"efbf0",-- -4161
x"eec30",-- -4413
x"ee370",-- -4553
x"edac0",-- -4692
x"ecff0",-- -4865
x"eda10",-- -4703
x"f0320",-- -4046
x"f3ef0",-- -3089
x"f87f0",-- -1921
x"fe260",-- -474
x"03f30",-- 1011
x"08200",-- 2080
x"0b4e0",-- 2894
x"0e250",-- 3621
x"0e750",-- 3701
x"0cd20",-- 3282
x"0a4a0",-- 2634
x"07f90",-- 2041
x"062b0",-- 1579
x"04e00",-- 1248
x"040d0",-- 1037
x"02fa0",-- 762
x"02d10",-- 721
x"036a0",-- 874
x"031a0",-- 794
x"018b0",-- 395
x"002b0",-- 43
x"fef50",-- -267
x"fe030",-- -509
x"fd970",-- -617
x"feaf0",-- -337
x"00e40",-- 228
x"039a0",-- 922
x"07850",-- 1925
x"0c050",-- 3077
x"11620",-- 4450
x"16b30",-- 5811
x"1b9c0",-- 7068
x"1fbf0",-- 8127
x"23740",-- 9076
x"277b0",-- 10107
x"2aab0",-- 10923
x"2b8f0",-- 11151
x"29eb0",-- 10731
x"267e0",-- 9854
x"22320",-- 8754
x"1cfc0",-- 7420
x"156f0",-- 5487
x"0ad70",-- 2775
x"fe500",-- -432
x"f1450",-- -3771
x"e53d0",-- -6851
x"dba00",-- -9312
x"d5d60",-- -10794
x"d1d40",-- -11820
x"ceda0",-- -12582
x"ced60",-- -12586
x"d36b0",-- -11413
x"da640",-- -9628
x"e0a60",-- -8026
x"e4990",-- -7015
x"e8080",-- -6136
x"ed4d0",-- -4787
x"f5470",-- -2745
x"fdef0",-- -529
x"05790",-- 1401
x"0d400",-- 3392
x"167c0",-- 5756
x"1f280",-- 7976
x"26200",-- 9760
x"2a470",-- 10823
x"2a270",-- 10791
x"24f10",-- 9457
x"1c0c0",-- 7180
x"116f0",-- 4463
x"05990",-- 1433
x"f9520",-- -1710
x"ed1a0",-- -4838
x"e1f70",-- -7689
x"dab90",-- -9543
x"d8280",-- -10200
x"d83f0",-- -10177
x"d9340",-- -9932
x"dad20",-- -9518
x"de080",-- -8696
x"e2800",-- -7552
x"e6690",-- -6551
x"ea4b0",-- -5557
x"edc90",-- -4663
x"f2120",-- -3566
x"f7ab0",-- -2133
x"fe7d0",-- -387
x"05d10",-- 1489
x"0d310",-- 3377
x"134f0",-- 4943
x"16320",-- 5682
x"17bc0",-- 6076
x"18a40",-- 6308
x"192b0",-- 6443
x"16ae0",-- 5806
x"11100",-- 4368
x"0b770",-- 2935
x"076a0",-- 1898
x"051c0",-- 1308
x"01060",-- 262
x"fbba0",-- -1094
x"f6ac0",-- -2388
x"f2e60",-- -3354
x"f0260",-- -4058
x"ed930",-- -4717
x"ece90",-- -4887
x"ede50",-- -4635
x"ef100",-- -4336
x"f1330",-- -3789
x"f60a0",-- -2550
x"fc750",-- -907
x"020a0",-- 522
x"04580",-- 1112
x"050b0",-- 1291
x"061e0",-- 1566
x"072b0",-- 1835
x"072b0",-- 1835
x"04200",-- 1056
x"01bd0",-- 445
x"01c40",-- 452
x"02f40",-- 756
x"03860",-- 902
x"03620",-- 866
x"030d0",-- 781
x"01ec0",-- 492
x"00200",-- 32
x"fe300",-- -464
x"fc3f0",-- -961
x"fa0f0",-- -1521
x"f86b0",-- -1941
x"f7a40",-- -2140
x"f9270",-- -1753
x"fcd70",-- -809
x"00960",-- 150
x"031a0",-- 794
x"04cc0",-- 1228
x"08050",-- 2053
x"0b620",-- 2914
x"0d2c0",-- 3372
x"0d8d0",-- 3469
x"0d270",-- 3367
x"0d380",-- 3384
x"0dd60",-- 3542
x"0f630",-- 3939
x"11a60",-- 4518
x"15380",-- 5432
x"191a0",-- 6426
x"1c130",-- 7187
x"1f320",-- 7986
x"21f30",-- 8691
x"263b0",-- 9787
x"278f0",-- 10127
x"248d0",-- 9357
x"1d6c0",-- 7532
x"16130",-- 5651
x"127d0",-- 4733
x"0bfe0",-- 3070
x"032c0",-- 812
x"f6910",-- -2415
x"ec0b0",-- -5109
x"e4a30",-- -7005
x"e04b0",-- -8117
x"def10",-- -8463
x"db9a0",-- -9318
x"dafa0",-- -9478
x"db8e0",-- -9330
x"def30",-- -8461
x"e3480",-- -7352
x"e8f30",-- -5901
x"ecca0",-- -4918
x"eda20",-- -4702
x"f1bb0",-- -3653
x"fa170",-- -1513
x"05090",-- 1289
x"0cd70",-- 3287
x"138d0",-- 5005
x"182c0",-- 6188
x"1cb10",-- 7345
x"1f690",-- 8041
x"1ce70",-- 7399
x"15910",-- 5521
x"0b040",-- 2820
x"01b00",-- 432
x"f7d50",-- -2091
x"ef310",-- -4303
x"e8e60",-- -5914
x"e4060",-- -7162
x"dfbf0",-- -8257
x"de4e0",-- -8626
x"e12c0",-- -7892
x"e4800",-- -7040
x"e7740",-- -6284
x"e9bb0",-- -5701
x"ed8e0",-- -4722
x"f3070",-- -3321
x"fa1e0",-- -1506
x"ff920",-- -110
x"02e60",-- 742
x"069d0",-- 1693
x"0a000",-- 2560
x"0ce60",-- 3302
x"0d830",-- 3459
x"0cbb0",-- 3259
x"0b060",-- 2822
x"06440",-- 1604
x"006b0",-- 107
x"fd920",-- -622
x"fe820",-- -382
x"007d0",-- 125
x"fdb20",-- -590
x"f8990",-- -1895
x"f7600",-- -2208
x"fa8e0",-- -1394
x"fc080",-- -1016
x"f8fc0",-- -1796
x"f56f0",-- -2705
x"f6ad0",-- -2387
x"fb4a0",-- -1206
x"fee40",-- -284
x"02b10",-- 689
x"05f40",-- 1524
x"09880",-- 2440
x"08320",-- 2098
x"06410",-- 1601
x"06930",-- 1683
x"05400",-- 1344
x"02170",-- 535
x"faeb0",-- -1301
x"f8080",-- -2040
x"f9700",-- -1680
x"fa760",-- -1418
x"f8ee0",-- -1810
x"f5790",-- -2695
x"f5770",-- -2697
x"f7e50",-- -2075
x"f84e0",-- -1970
x"f8190",-- -2023
x"f95b0",-- -1701
x"fb850",-- -1147
x"fdcc0",-- -564
x"ff630",-- -157
x"03da0",-- 986
x"072b0",-- 1835
x"07ec0",-- 2028
x"074c0",-- 1868
x"070b0",-- 1803
x"09f60",-- 2550
x"0aa70",-- 2727
x"08d60",-- 2262
x"06b60",-- 1718
x"078a0",-- 1930
x"0a460",-- 2630
x"0ad60",-- 2774
x"096f0",-- 2415
x"08110",-- 2065
x"06e00",-- 1760
x"054e0",-- 1358
x"05150",-- 1301
x"06b80",-- 1720
x"0c460",-- 3142
x"134a0",-- 4938
x"1a1b0",-- 6683
x"21140",-- 8468
x"26520",-- 9810
x"2ad80",-- 10968
x"293f0",-- 10559
x"24c90",-- 9417
x"1dec0",-- 7660
x"18af0",-- 6319
x"173c0",-- 5948
x"100c0",-- 4108
x"06440",-- 1604
x"f9d10",-- -1583
x"f23e0",-- -3522
x"eb7c0",-- -5252
x"e2cd0",-- -7475
x"dc290",-- -9175
x"d8510",-- -10159
x"d9ac0",-- -9812
x"ddca0",-- -8758
x"e3d10",-- -7215
x"e9480",-- -5816
x"ee9d0",-- -4451
x"f1f10",-- -3599
x"f55e0",-- -2722
x"f9540",-- -1708
x"02030",-- 515
x"09d50",-- 2517
x"0e3e0",-- 3646
x"13850",-- 4997
x"18810",-- 6273
x"1cf60",-- 7414
x"1aa00",-- 6816
x"13bf0",-- 5055
x"0a1c0",-- 2588
x"00000",-- 0
x"f68c0",-- -2420
x"ed720",-- -4750
x"e5ac0",-- -6740
x"e0bc0",-- -8004
x"de140",-- -8684
x"dc5f0",-- -9121
x"dce70",-- -8985
x"dfde0",-- -8226
x"e4150",-- -7147
x"e6960",-- -6506
x"eb110",-- -5359
x"f2010",-- -3583
x"fa210",-- -1503
x"01dd0",-- 477
x"06e30",-- 1763
x"0afe0",-- 2814
x"0e0f0",-- 3599
x"0f8d0",-- 3981
x"0eb90",-- 3769
x"0be20",-- 3042
x"08db0",-- 2267
x"05830",-- 1411
x"02c00",-- 704
x"00690",-- 105
x"ff3f0",-- -193
x"fb9f0",-- -1121
x"f6260",-- -2522
x"f4d50",-- -2859
x"f7720",-- -2190
x"fb390",-- -1223
x"fafc0",-- -1284
x"f9630",-- -1693
x"f9330",-- -1741
x"fe890",-- -375
x"04be0",-- 1214
x"05d60",-- 1494
x"03810",-- 897
x"02d90",-- 729
x"075b0",-- 1883
x"09db0",-- 2523
x"0a2d0",-- 2605
x"07b00",-- 1968
x"04780",-- 1144
x"00440",-- 68
x"fd8f0",-- -625
x"fd670",-- -665
x"fb480",-- -1208
x"f9200",-- -1760
x"f6a30",-- -2397
x"f62b0",-- -2517
x"f8890",-- -1911
x"faf20",-- -1294
x"fa320",-- -1486
x"f7c60",-- -2106
x"f8030",-- -2045
x"fb180",-- -1256
x"fdd60",-- -554
x"fef00",-- -272
x"00960",-- 150
x"02640",-- 612
x"04340",-- 1076
x"05ce0",-- 1486
x"05fe0",-- 1534
x"04140",-- 1044
x"01fd0",-- 509
x"01260",-- 294
x"018d0",-- 397
x"04250",-- 1061
x"068b0",-- 1675
x"06d90",-- 1753
x"06f70",-- 1783
x"08a70",-- 2215
x"09f80",-- 2552
x"08c20",-- 2242
x"06d10",-- 1745
x"05b70",-- 1463
x"08c30",-- 2243
x"109b0",-- 4251
x"19030",-- 6403
x"213c0",-- 8508
x"26e00",-- 9952
x"2a6f0",-- 10863
x"2b050",-- 11013
x"29300",-- 10544
x"25bf0",-- 9663
x"1d230",-- 7459
x"149d0",-- 5277
x"0f330",-- 3891
x"0c070",-- 3079
x"04ef0",-- 1263
x"f9950",-- -1643
x"ede50",-- -4635
x"e2260",-- -7642
x"db4f0",-- -9393
x"d8f30",-- -9997
x"d9ac0",-- -9812
x"dbe50",-- -9243
x"e1320",-- -7886
x"e83c0",-- -6084
x"efa60",-- -4186
x"f6850",-- -2427
x"fa2a0",-- -1494
x"fb2e0",-- -1234
x"fcbb0",-- -837
x"03ec0",-- 1004
x"0d8d0",-- 3469
x"16630",-- 5731
x"1b320",-- 6962
x"1d140",-- 7444
x"1b4b0",-- 6987
x"15ab0",-- 5547
x"0d720",-- 3442
x"01c70",-- 455
x"f5700",-- -2704
x"ea5f0",-- -5537
x"e2d30",-- -7469
x"dec40",-- -8508
x"dddb0",-- -8741
x"dc3f0",-- -9153
x"da4b0",-- -9653
x"da280",-- -9688
x"dd280",-- -8920
x"e2cd0",-- -7475
x"e9680",-- -5784
x"f1360",-- -3786
x"fa5a0",-- -1446
x"04b40",-- 1204
x"0cff0",-- 3327
x"12770",-- 4727
x"13ba0",-- 5050
x"11ff0",-- 4607
x"0eb40",-- 3764
x"0acf0",-- 2767
x"07a60",-- 1958
x"05530",-- 1363
x"02690",-- 617
x"fed40",-- -300
x"fbe00",-- -1056
x"f9c40",-- -1596
x"f7680",-- -2200
x"f2f20",-- -3342
x"ee670",-- -4505
x"eb520",-- -5294
x"f09b0",-- -3941
x"f7f90",-- -2055
x"fff40",-- -12
x"04350",-- 1077
x"07cb0",-- 1995
x"08910",-- 2193
x"04260",-- 1062
x"07940",-- 1940
x"08910",-- 2193
x"0bc70",-- 3015
x"069f0",-- 1695
x"073b0",-- 1851
x"0c570",-- 3159
x"0b810",-- 2945
x"09b70",-- 2487
x"fd400",-- -704
x"f7750",-- -2187
x"f3b80",-- -3144
x"f3ac0",-- -3156
x"f5040",-- -2812
x"f5100",-- -2800
x"f9db0",-- -1573
x"faee0",-- -1298
x"f97e0",-- -1666
x"fab60",-- -1354
x"fae40",-- -1308
x"f9fd0",-- -1539
x"f8b90",-- -1863
x"fb1b0",-- -1253
x"02990",-- 665
x"070b0",-- 1803
x"096a0",-- 2410
x"07920",-- 1938
x"05fe0",-- 1534
x"05490",-- 1353
x"02e00",-- 736
x"ffd10",-- -47
x"ff360",-- -202
x"025c0",-- 604
x"05580",-- 1368
x"086d0",-- 2157
x"0b580",-- 2904
x"0d970",-- 3479
x"0a230",-- 2595
x"06be0",-- 1726
x"047d0",-- 1149
x"06390",-- 1593
x"0c5e0",-- 3166
x"12a70",-- 4775
x"198a0",-- 6538
x"1f800",-- 8064
x"27790",-- 10105
x"2bd40",-- 11220
x"2bb70",-- 11191
x"273c0",-- 10044
x"213c0",-- 8508
x"1a6b0",-- 6763
x"15cb0",-- 5579
x"133b0",-- 4923
x"0c870",-- 3207
x"018a0",-- 394
x"f2b40",-- -3404
x"e71b0",-- -6373
x"dd3c0",-- -8900
x"d81f0",-- -10209
x"d7aa0",-- -10326
x"db570",-- -9385
x"e2920",-- -7534
x"e8a00",-- -5984
x"ef1f0",-- -4321
x"f4580",-- -2984
x"f7950",-- -2155
x"f8780",-- -1928
x"f97e0",-- -1666
x"fee40",-- -284
x"09cc0",-- 2508
x"14310",-- 5169
x"1bab0",-- 7083
x"1e960",-- 7830
x"1c7c0",-- 7292
x"16720",-- 5746
x"0c500",-- 3152
x"01650",-- 357
x"f6de0",-- -2338
x"eeaf0",-- -4433
x"e7de0",-- -6178
x"e2e70",-- -7449
x"e0830",-- -8061
x"dd6e0",-- -8850
x"d9d70",-- -9769
x"d6f00",-- -10512
x"d7640",-- -10396
x"dd4f0",-- -8881
x"e5f40",-- -6668
x"f1010",-- -3839
x"fcf80",-- -776
x"077b0",-- 1915
x"0f510",-- 3921
x"13360",-- 4918
x"134a0",-- 4938
x"10f70",-- 4343
x"0db20",-- 3506
x"0a200",-- 2592
x"07e70",-- 2023
x"06d90",-- 1753
x"04930",-- 1171
x"001c0",-- 28
x"faf20",-- -1294
x"f52f0",-- -2769
x"f0d70",-- -3881
x"edfc0",-- -4612
x"ed4d0",-- -4787
x"eeb40",-- -4428
x"ee670",-- -4505
x"f36a0",-- -3222
x"fd4e0",-- -690
x"08660",-- 2150
x"0b620",-- 2914
x"0b5e0",-- 2910
x"07590",-- 1881
x"05420",-- 1346
x"0be90",-- 3049
x"0ed20",-- 3794
x"10a90",-- 4265
x"09720",-- 2418
x"0a080",-- 2568
x"0ad70",-- 2775
x"08350",-- 2101
x"040d0",-- 1037
x"f8350",-- -1995
x"f1f90",-- -3591
x"ee080",-- -4600
x"f2430",-- -3517
x"f7df0",-- -2081
x"f78d0",-- -2163
x"f92c0",-- -1748
x"f6ff0",-- -2305
x"f6730",-- -2445
x"f9830",-- -1661
x"f9310",-- -1743
x"fa3f0",-- -1473
x"fb7b0",-- -1157
x"01ee0",-- 494
x"08870",-- 2183
x"0ae00",-- 2784
x"0ac80",-- 2760
x"06cc0",-- 1740
x"037e0",-- 894
x"01620",-- 354
x"00940",-- 148
x"00750",-- 117
x"00b60",-- 182
x"02ad0",-- 685
x"05b30",-- 1459
x"080f0",-- 2063
x"09a90",-- 2473
x"08580",-- 2136
x"06900",-- 1680
x"07900",-- 1936
x"0aaa0",-- 2730
x"0d330",-- 3379
x"11060",-- 4358
x"14b90",-- 5305
x"185a0",-- 6234
x"1d690",-- 7529
x"22950",-- 8853
x"28330",-- 10291
x"2a060",-- 10758
x"29650",-- 10597
x"253a0",-- 9530
x"1ec50",-- 7877
x"19e10",-- 6625
x"13bf0",-- 5055
x"07470",-- 1863
x"f6870",-- -2425
x"e9600",-- -5792
x"e2c30",-- -7485
x"dfab0",-- -8277
x"df750",-- -8331
x"e0a10",-- -8031
x"e1630",-- -7837
x"e5770",-- -6793
x"e9ec0",-- -5652
x"ee6b0",-- -4501
x"f1a10",-- -3679
x"f4b60",-- -2890
x"f88c0",-- -1908
x"fe8a0",-- -374
x"08d70",-- 2263
x"11f50",-- 4597
x"16820",-- 5762
x"16b60",-- 5814
x"15760",-- 5494
x"12690",-- 4713
x"0d3a0",-- 3386
x"06b40",-- 1716
x"ffd00",-- -48
x"f88c0",-- -1908
x"f1f40",-- -3596
x"eab70",-- -5449
x"e31d0",-- -7395
x"dd130",-- -8941
x"d7950",-- -10347
x"d4b50",-- -11083
x"d6500",-- -10672
x"dd1e0",-- -8930
x"e6170",-- -6633
x"ef8d0",-- -4211
x"f8d90",-- -1831
x"00f00",-- 240
x"08020",-- 2050
x"0c410",-- 3137
x"0e200",-- 3616
x"0e9b0",-- 3739
x"0e700",-- 3696
x"0d9f0",-- 3487
x"0b970",-- 2967
x"089d0",-- 2205
x"04280",-- 1064
x"fe6e0",-- -402
x"f8480",-- -1976
x"f3920",-- -3182
x"f0e30",-- -3869
x"efea0",-- -4118
x"f0960",-- -3946
x"f33d0",-- -3267
x"f6350",-- -2507
x"f9e70",-- -1561
x"f8930",-- -1901
x"f9010",-- -1791
x"00020",-- 2
x"08d10",-- 2257
x"0fd20",-- 4050
x"09740",-- 2420
x"09770",-- 2423
x"0d310",-- 3377
x"11620",-- 4450
x"10140",-- 4116
x"05860",-- 1414
x"038f0",-- 911
x"00730",-- 115
x"01120",-- 274
x"00960",-- 150
x"fb9a0",-- -1126
x"f8140",-- -2028
x"f19c0",-- -3684
x"ef740",-- -4236
x"f3b50",-- -3147
x"f54f0",-- -2737
x"f6b70",-- -2377
x"f48c0",-- -2932
x"f7560",-- -2218
x"ff010",-- -255
x"00550",-- 85
x"00700",-- 112
x"fd9c0",-- -612
x"ffd50",-- -43
x"03510",-- 849
x"04dc0",-- 1244
x"06760",-- 1654
x"06280",-- 1576
x"05d60",-- 1494
x"04940",-- 1172
x"03740",-- 884
x"03d50",-- 981
x"031f0",-- 799
x"00800",-- 128
x"00bc0",-- 188
x"03ec0",-- 1004
x"09030",-- 2307
x"0b170",-- 2839
x"0a7f0",-- 2687
x"0b4f0",-- 2895
x"0d920",-- 3474
x"0f0d0",-- 3853
x"105e0",-- 4190
x"136c0",-- 4972
x"198a0",-- 6538
x"207e0",-- 8318
x"24d80",-- 9432
x"29870",-- 10631
x"2b410",-- 11073
x"29fa0",-- 10746
x"21dc0",-- 8668
x"174c0",-- 5964
x"116c0",-- 4460
x"09030",-- 2307
x"fd4c0",-- -692
x"ed070",-- -4857
x"e3cf0",-- -7217
x"e1cc0",-- -7732
x"e0ce0",-- -7986
x"e1cc0",-- -7732
x"e2120",-- -7662
x"e56a0",-- -6806
x"e8290",-- -6103
x"ebc70",-- -5177
x"f1200",-- -3808
x"f69e0",-- -2402
x"fb590",-- -1191
x"ffbf0",-- -65
x"05c60",-- 1478
x"0de50",-- 3557
x"13ce0",-- 5070
x"146b0",-- 5227
x"11c10",-- 4545
x"0e280",-- 3624
x"0be20",-- 3042
x"06c20",-- 1730
x"01100",-- 272
x"fade0",-- -1314
x"f4140",-- -3052
x"ecc50",-- -4923
x"e4640",-- -7068
x"de870",-- -8569
x"da4e0",-- -9650
x"d7fc0",-- -10244
x"d88f0",-- -10097
x"ddea0",-- -8726
x"e69b0",-- -6501
x"f08e0",-- -3954
x"f86b0",-- -1941
x"ff2e0",-- -210
x"05560",-- 1366
x"0a7f0",-- 2687
x"0d7e0",-- 3454
x"0e0f0",-- 3599
x"0e520",-- 3666
x"0cb80",-- 3256
x"0ad70",-- 2775
x"06f90",-- 1785
x"02550",-- 597
x"fced0",-- -787
x"f7560",-- -2218
x"f30c0",-- -3316
x"f0670",-- -3993
x"f1250",-- -3803
x"f2840",-- -3452
x"f5a40",-- -2652
x"f72f0",-- -2257
x"f61c0",-- -2532
x"f8980",-- -1896
x"000c0",-- 12
x"07860",-- 1926
x"0c690",-- 3177
x"0a980",-- 2712
x"08840",-- 2180
x"0c310",-- 3121
x"0de90",-- 3561
x"104d0",-- 4173
x"08a20",-- 2210
x"051c0",-- 1308
x"040f0",-- 1039
x"02430",-- 579
x"03010",-- 769
x"fc7b0",-- -901
x"f84b0",-- -1973
x"f23a0",-- -3526
x"f0bb0",-- -3909
x"f4fa0",-- -2822
x"f6490",-- -2487
x"f70b0",-- -2293
x"f7660",-- -2202
x"f7ab0",-- -2133
x"fc820",-- -894
x"fe030",-- -509
x"fd850",-- -635
x"fd540",-- -684
x"fe2a0",-- -470
x"03530",-- 851
x"05860",-- 1414
x"06960",-- 1686
x"05010",-- 1281
x"02030",-- 515
x"00ac0",-- 172
x"008e0",-- 142
x"01310",-- 305
x"01630",-- 355
x"00800",-- 128
x"018d0",-- 397
x"04580",-- 1112
x"06b60",-- 1718
x"08f20",-- 2290
x"07fd0",-- 2045
x"08820",-- 2178
x"0bfe0",-- 3070
x"0fc10",-- 4033
x"12cc0",-- 4812
x"13b90",-- 5049
x"15f30",-- 5619
x"18d10",-- 6353
x"1ddc0",-- 7644
x"23470",-- 9031
x"25ec0",-- 9708
x"28ba0",-- 10426
x"28830",-- 10371
x"24ab0",-- 9387
x"1afe0",-- 6910
x"122f0",-- 4655
x"08fa0",-- 2298
x"fc5c0",-- -932
x"ee490",-- -4535
x"e34f0",-- -7345
x"e0100",-- -8176
x"e21f0",-- -7649
x"e5c50",-- -6715
x"e5fb0",-- -6661
x"e8ed0",-- -5907
x"eb630",-- -5277
x"ee6b0",-- -4501
x"f0930",-- -3949
x"f5db0",-- -2597
x"fc190",-- -999
x"00160",-- 22
x"060f0",-- 1551
x"0c9a0",-- 3226
x"12770",-- 4727
x"11da0",-- 4570
x"0df80",-- 3576
x"08b40",-- 2228
x"05d60",-- 1494
x"02c50",-- 709
x"ff240",-- -220
x"fa110",-- -1519
x"f50c0",-- -2804
x"eeaf0",-- -4433
x"e63f0",-- -6593
x"e03d0",-- -8131
x"db410",-- -9407
x"da380",-- -9672
x"db250",-- -9435
x"e19a0",-- -7782
x"eabb0",-- -5445
x"f4460",-- -3002
x"fb600",-- -1184
x"00870",-- 135
x"05720",-- 1394
x"08a70",-- 2215
x"0b220",-- 2850
x"0ba60",-- 2982
x"0bd00",-- 3024
x"0b1d0",-- 2845
x"08af0",-- 2223
x"04230",-- 1059
x"ff240",-- -220
x"f9e70",-- -1561
x"f4bc0",-- -2884
x"f1700",-- -3728
x"f14c0",-- -3764
x"f3950",-- -3179
x"f6480",-- -2488
x"f98b0",-- -1653
x"fae60",-- -1306
x"f9040",-- -1788
x"fce10",-- -799
x"02ff0",-- 767
x"06f90",-- 1785
x"09e40",-- 2532
x"0afc0",-- 2812
x"10340",-- 4148
x"0f2c0",-- 3884
x"0d7c0",-- 3452
x"0a340",-- 2612
x"03830",-- 899
x"026b0",-- 619
x"ff580",-- -168
x"ff2e0",-- -210
x"fd970",-- -617
x"fa480",-- -1464
x"f7fb0",-- -2053
x"f48a0",-- -2934
x"f4e90",-- -2839
x"f5ef0",-- -2577
x"f4700",-- -2960
x"f6d40",-- -2348
x"f9f10",-- -1551
x"fd680",-- -664
x"00000",-- 0
x"ffa10",-- -95
x"006b0",-- 107
x"ff7c0",-- -132
x"00610",-- 97
x"01620",-- 354
x"01df0",-- 479
x"028a0",-- 650
x"02350",-- 565
x"02260",-- 550
x"02390",-- 569
x"01bf0",-- 447
x"005a0",-- 90
x"00610",-- 97
x"00e90",-- 233
x"03310",-- 817
x"045c0",-- 1116
x"06610",-- 1633
x"09330",-- 2355
x"0b6c0",-- 2924
x"0df80",-- 3576
x"0fe10",-- 4065
x"10cc0",-- 4300
x"11260",-- 4390
x"13d30",-- 5075
x"17d20",-- 6098
x"1cd30",-- 7379
x"20e80",-- 8424
x"243b0",-- 9275
x"25dc0",-- 9692
x"26b10",-- 9905
x"244c0",-- 9292
x"1cd10",-- 7377
x"15790",-- 5497
x"0eac0",-- 3756
x"064e0",-- 1614
x"fb420",-- -1214
x"ef700",-- -4240
x"e7660",-- -6298
x"e2c90",-- -7479
x"e3930",-- -7277
x"e6f70",-- -6409
x"e9040",-- -5884
x"ec0f0",-- -5105
x"ee7a0",-- -4486
x"f2530",-- -3501
x"f64e0",-- -2482
x"fa4e0",-- -1458
x"fc9e0",-- -866
x"fe9d0",-- -355
x"03e40",-- 996
x"09bc0",-- 2492
x"0c720",-- 3186
x"0b920",-- 2962
x"08930",-- 2195
x"04500",-- 1104
x"00930",-- 147
x"fd0e0",-- -754
x"f98d0",-- -1651
x"f5090",-- -2807
x"f07f0",-- -3969
x"ebf10",-- -5135
x"e7840",-- -6268
x"e38e0",-- -7282
x"e0550",-- -8107
x"df4a0",-- -8374
x"e1770",-- -7817
x"e8170",-- -6121
x"efe80",-- -4120
x"f7830",-- -2173
x"fe3f0",-- -449
x"03850",-- 901
x"06d10",-- 1745
x"08aa0",-- 2218
x"0a0a0",-- 2570
x"096a0",-- 2410
x"07c90",-- 1993
x"05400",-- 1344
x"02800",-- 640
x"feaf0",-- -337
x"f9e90",-- -1559
x"f57a0",-- -2694
x"f32a0",-- -3286
x"f3470",-- -3257
x"f4a70",-- -2905
x"f6780",-- -2440
x"f8bc0",-- -1860
x"fc980",-- -872
x"003f0",-- 63
x"038d0",-- 909
x"06210",-- 1569
x"08cd0",-- 2253
x"09ee0",-- 2542
x"0bb00",-- 2992
x"0c220",-- 3106
x"0c610",-- 3169
x"0b210",-- 2849
x"08530",-- 2131
x"05cc0",-- 1484
x"023f0",-- 575
x"008a0",-- 138
x"fd790",-- -647
x"fabc0",-- -1348
x"f8c10",-- -1855
x"f76b0",-- -2197
x"f69e0",-- -2402
x"f68c0",-- -2420
x"f6c80",-- -2360
x"f89d0",-- -1891
x"f9700",-- -1680
x"fb0c0",-- -1268
x"fd1a0",-- -742
x"fe250",-- -475
x"00280",-- 40
x"008c0",-- 140
x"018d0",-- 397
x"02350",-- 565
x"025d0",-- 605
x"01ba0",-- 442
x"00f70",-- 247
x"01350",-- 309
x"01d60",-- 470
x"01030",-- 259
x"00d20",-- 210
x"008f0",-- 143
x"01310",-- 305
x"02750",-- 629
x"02ef0",-- 751
x"04820",-- 1154
x"05bd0",-- 1469
x"08be0",-- 2238
x"0bb00",-- 2992
x"0e900",-- 3728
x"11c90",-- 4553
x"14570",-- 5207
x"145c0",-- 5212
x"14730",-- 5235
x"146e0",-- 5230
x"19650",-- 6501
x"1dd30",-- 7635
x"21aa0",-- 8618
x"24b50",-- 9397
x"23460",-- 9030
x"220a0",-- 8714
x"19960",-- 6550
x"13df0",-- 5087
x"0e5e0",-- 3678
x"07a30",-- 1955
x"fd8b0",-- -629
x"f1ab0",-- -3669
x"eaee0",-- -5394
x"e7e00",-- -6176
x"e8030",-- -6141
x"e60b0",-- -6645
x"e7b60",-- -6218
x"eb9d0",-- -5219
x"f1c50",-- -3643
x"f54d0",-- -2739
x"f8d50",-- -1835
x"fc120",-- -1006
x"fca70",-- -857
x"fe4e0",-- -434
x"00260",-- 38
x"05440",-- 1348
x"06e60",-- 1766
x"069a0",-- 1690
x"045a0",-- 1114
x"02c00",-- 704
x"ff9a0",-- -102
x"fa430",-- -1469
x"f5c00",-- -2624
x"f1740",-- -3724
x"f00b0",-- -4085
x"ed0e0",-- -4850
x"ea4b0",-- -5557
x"e7650",-- -6299
x"e5600",-- -6816
x"e4170",-- -7145
x"e5840",-- -6780
x"ea670",-- -5529
x"f0100",-- -4080
x"f6f50",-- -2315
x"fc8a0",-- -886
x"031f0",-- 799
x"07950",-- 1941
x"09800",-- 2432
x"08080",-- 2056
x"05b80",-- 1464
x"03330",-- 819
x"00a70",-- 167
x"ff7e0",-- -130
x"fd470",-- -697
x"fabe0",-- -1346
x"f6be0",-- -2370
x"f3c00",-- -3136
x"f31a0",-- -3302
x"f5840",-- -2684
x"f7660",-- -2202
x"fa7d0",-- -1411
x"fe030",-- -509
x"02120",-- 530
x"06910",-- 1681
x"09420",-- 2370
x"0a210",-- 2593
x"0a0d0",-- 2573
x"09540",-- 2388
x"0a1c0",-- 2588
x"0a820",-- 2690
x"09e00",-- 2528
x"08440",-- 2116
x"03e90",-- 1001
x"022b0",-- 555
x"fde50",-- -539
x"fb7b0",-- -1157
x"f8d20",-- -1838
x"f7020",-- -2302
x"f79c0",-- -2148
x"f7b20",-- -2126
x"f88c0",-- -1908
x"f97c0",-- -1668
x"f98b0",-- -1653
x"fa0c0",-- -1524
x"fbb20",-- -1102
x"fce60",-- -794
x"ffb80",-- -72
x"001e0",-- 30
x"019f0",-- 415
x"02350",-- 565
x"02c80",-- 712
x"02800",-- 640
x"002a0",-- 42
x"ff9c0",-- -100
x"ff110",-- -239
x"ffe90",-- -23
x"00c10",-- 193
x"020f0",-- 527
x"02de0",-- 734
x"03bf0",-- 959
x"03ea0",-- 1002
x"04b10",-- 1201
x"061b0",-- 1563
x"07a10",-- 1953
x"0a630",-- 2659
x"0d470",-- 3399
x"10a20",-- 4258
x"14050",-- 5125
x"148b0",-- 5259
x"14050",-- 5125
x"133f0",-- 4927
x"15120",-- 5394
x"19690",-- 6505
x"1e700",-- 7792
x"233d0",-- 9021
x"23c40",-- 9156
x"21d00",-- 8656
x"1ce00",-- 7392
x"16c20",-- 5826
x"12640",-- 4708
x"0ae50",-- 2789
x"fee10",-- -287
x"f1200",-- -3808
x"ecfa0",-- -4870
x"eced0",-- -4883
x"ea780",-- -5512
x"e6a80",-- -6488
x"e6f50",-- -6411
x"ec6a0",-- -5014
x"f16d0",-- -3731
x"f54a0",-- -2742
x"f6750",-- -2443
x"f9130",-- -1773
x"fad20",-- -1326
x"ff180",-- -232
x"01d10",-- 465
x"05630",-- 1379
x"053d0",-- 1341
x"036f0",-- 879
x"030e0",-- 782
x"023e0",-- 574
x"ff970",-- -105
x"f8930",-- -1901
x"f4a70",-- -2905
x"f2a50",-- -3419
x"f23f0",-- -3521
x"ef250",-- -4315
x"eb240",-- -5340
x"e7830",-- -6269
x"e5d60",-- -6698
x"e61c0",-- -6628
x"e6b00",-- -6480
x"ea0d0",-- -5619
x"ef450",-- -4283
x"f6460",-- -2490
x"fcc50",-- -827
x"02840",-- 644
x"069a0",-- 1690
x"06ff0",-- 1791
x"05260",-- 1318
x"04250",-- 1061
x"04260",-- 1062
x"03450",-- 837
x"00640",-- 100
x"fe050",-- -507
x"fbc40",-- -1084
x"f9330",-- -1741
x"f4e60",-- -2842
x"f2340",-- -3532
x"f2730",-- -3469
x"f56b0",-- -2709
x"f9270",-- -1753
x"fd060",-- -762
x"02c00",-- 704
x"06d20",-- 1746
x"09130",-- 2323
x"09770",-- 2423
x"0a030",-- 2563
x"0a4f0",-- 2639
x"0b040",-- 2820
x"0a3c0",-- 2620
x"0a4a0",-- 2634
x"08db0",-- 2267
x"069d0",-- 1693
x"039a0",-- 922
x"fe410",-- -447
x"fbae0",-- -1106
x"f8350",-- -1995
x"f6c00",-- -2368
x"f6850",-- -2427
x"f7750",-- -2187
x"f9090",-- -1783
x"f9b00",-- -1616
x"fa1b0",-- -1509
x"fa6b0",-- -1429
x"fa7d0",-- -1411
x"fbd30",-- -1069
x"fe300",-- -464
x"00110",-- 17
x"02b10",-- 689
x"03920",-- 914
x"037c0",-- 892
x"028f0",-- 655
x"01510",-- 337
x"009d0",-- 157
x"ffa60",-- -90
x"ff310",-- -207
x"fff60",-- -10
x"01c70",-- 455
x"02aa0",-- 682
x"03120",-- 786
x"02aa0",-- 682
x"03450",-- 837
x"04b90",-- 1209
x"07090",-- 1801
x"0a540",-- 2644
x"0dc60",-- 3526
x"112b0",-- 4395
x"13650",-- 4965
x"14310",-- 5169
x"12280",-- 4648
x"124d0",-- 4685
x"12c00",-- 4800
x"17600",-- 5984
x"1c570",-- 7255
x"21d20",-- 8658
x"255a0",-- 9562
x"22400",-- 8768
x"1e390",-- 7737
x"16950",-- 5781
x"11310",-- 4401
x"0a980",-- 2712
x"02710",-- 625
x"f7a80",-- -2136
x"eeb70",-- -4425
x"ed0e0",-- -4850
x"ed3b0",-- -4805
x"eb3b0",-- -5317
x"e8780",-- -6024
x"e9ae0",-- -5714
x"ec7d0",-- -4995
x"f2750",-- -3467
x"f7270",-- -2265
x"fb5e0",-- -1186
x"fc080",-- -1016
x"fc070",-- -1017
x"ff650",-- -155
x"02b10",-- 689
x"03fe0",-- 1022
x"01080",-- 264
x"ff670",-- -153
x"ff580",-- -168
x"ff400",-- -192
x"fc4d0",-- -947
x"f7070",-- -2297
x"f30b0",-- -3317
x"f0bb0",-- -3909
x"eef70",-- -4361
x"ec870",-- -4985
x"ea870",-- -5497
x"e8170",-- -6121
x"e7450",-- -6331
x"e8d40",-- -5932
x"ec560",-- -5034
x"efbf0",-- -4161
x"f3a40",-- -3164
x"f8dc0",-- -1828
x"ff2b0",-- -213
x"04dc0",-- 1244
x"064b0",-- 1611
x"057c0",-- 1404
x"04340",-- 1076
x"045d0",-- 1117
x"03880",-- 904
x"ffdf0",-- -33
x"fcb40",-- -844
x"fa5f0",-- -1441
x"f8df0",-- -1825
x"f6840",-- -2428
x"f4eb0",-- -2837
x"f5380",-- -2760
x"f6820",-- -2430
x"f9860",-- -1658
x"fcff0",-- -769
x"00e10",-- 225
x"049d0",-- 1181
x"07710",-- 1905
x"08a50",-- 2213
x"0a4d0",-- 2637
x"0bd00",-- 3024
x"0c030",-- 3075
x"0ae10",-- 2785
x"09490",-- 2377
x"07f60",-- 2038
x"058d0",-- 1421
x"02ea0",-- 746
x"ff710",-- -143
x"fc730",-- -909
x"fa000",-- -1536
x"f9330",-- -1741
x"f8fc0",-- -1796
x"f8ac0",-- -1876
x"f8fd0",-- -1795
x"f8e10",-- -1823
x"f9e40",-- -1564
x"fb0b0",-- -1269
x"fc1e0",-- -994
x"fd020",-- -766
x"fddd0",-- -547
x"000c0",-- 12
x"01dd0",-- 477
x"028a0",-- 650
x"028f0",-- 655
x"01800",-- 384
x"01360",-- 310
x"013b0",-- 315
x"00d20",-- 210
x"00bc0",-- 188
x"006c0",-- 108
x"01490",-- 329
x"02b10",-- 689
x"03880",-- 904
x"03fb0",-- 1019
x"038b0",-- 907
x"04c20",-- 1218
x"07a60",-- 1958
x"0b120",-- 2834
x"0e4a0",-- 3658
x"10390",-- 4153
x"12d60",-- 4822
x"13820",-- 4994
x"134f0",-- 4943
x"12180",-- 4632
x"136f0",-- 4975
x"15e40",-- 5604
x"19b70",-- 6583
x"1efc0",-- 7932
x"240c0",-- 9228
x"242a0",-- 9258
x"1fb20",-- 8114
x"18050",-- 6149
x"12ac0",-- 4780
x"0e5c0",-- 3676
x"03db0",-- 987
x"f78d0",-- -2163
x"ecda0",-- -4902
x"ec9e0",-- -4962
x"ec150",-- -5099
x"eb9c0",-- -5220
x"e9970",-- -5737
x"eb7c0",-- -5252
x"ef3b0",-- -4293
x"f39d0",-- -3171
x"f78d0",-- -2163
x"f9970",-- -1641
x"fb310",-- -1231
x"fc390",-- -967
x"01310",-- 305
x"03990",-- 921
x"04cc0",-- 1228
x"01420",-- 322
x"ff4e0",-- -178
x"feda0",-- -294
x"fd330",-- -717
x"f9650",-- -1691
x"f4550",-- -2987
x"f2780",-- -3464
x"f1450",-- -3771
x"f0be0",-- -3906
x"ed700",-- -4752
x"ea5b0",-- -5541
x"e8150",-- -6123
x"e86a0",-- -6038
x"e9ea0",-- -5654
x"eceb0",-- -4885
x"f0d70",-- -3881
x"f56f0",-- -2705
x"fb2f0",-- -1233
x"00fc0",-- 252
x"04b40",-- 1204
x"045c0",-- 1116
x"038d0",-- 909
x"033b0",-- 827
x"045a0",-- 1114
x"02e00",-- 736
x"fff10",-- -15
x"fd400",-- -704
x"fb450",-- -1211
x"f9860",-- -1658
x"f5ef0",-- -2577
x"f3b30",-- -3149
x"f3900",-- -3184
x"f6070",-- -2553
x"f9c90",-- -1591
x"fe350",-- -459
x"03220",-- 802
x"06200",-- 1568
x"086b0",-- 2155
x"09ee0",-- 2542
x"0a980",-- 2712
x"0b760",-- 2934
x"0af00",-- 2800
x"0a4a0",-- 2634
x"0a660",-- 2662
x"096c0",-- 2412
x"06bd0",-- 1725
x"02750",-- 629
x"fda40",-- -604
x"fb880",-- -1144
x"f97f0",-- -1665
x"f8a50",-- -1883
x"f8170",-- -2025
x"f8730",-- -1933
x"fa3c0",-- -1476
x"fac00",-- -1344
x"fb560",-- -1194
x"fb620",-- -1182
x"fb760",-- -1162
x"fc750",-- -907
x"fdf90",-- -519
x"ffb20",-- -78
x"02730",-- 627
x"02f70",-- 759
x"03330",-- 819
x"028f0",-- 655
x"020d0",-- 525
x"01540",-- 340
x"003f0",-- 63
x"00440",-- 68
x"003c0",-- 60
x"004e0",-- 78
x"00800",-- 128
x"012e0",-- 302
x"01530",-- 339
x"02c10",-- 705
x"03fb0",-- 1019
x"06b60",-- 1718
x"09740",-- 2420
x"0ce80",-- 3304
x"0fd30",-- 4051
x"12180",-- 4632
x"14360",-- 5174
x"136a0",-- 4970
x"11e70",-- 4583
x"10e00",-- 4320
x"132c0",-- 4908
x"17d20",-- 6098
x"1d2b0",-- 7467
x"219b0",-- 8603
x"224b0",-- 8779
x"1fdf0",-- 8159
x"1c390",-- 7225
x"14eb0",-- 5355
x"0eac0",-- 3756
x"07590",-- 1881
x"ff8d0",-- -115
x"f4b20",-- -2894
x"eddb0",-- -4645
x"ed900",-- -4720
x"edc90",-- -4663
x"ecfa0",-- -4870
x"ea290",-- -5591
x"ed330",-- -4813
x"f1c20",-- -3646
x"f80c0",-- -2036
x"f9bc0",-- -1604
x"fbb20",-- -1102
x"fc200",-- -992
x"ff440",-- -188
x"02430",-- 579
x"01d00",-- 464
x"00500",-- 80
x"fdf60",-- -522
x"fe2d0",-- -467
x"fc4d0",-- -947
x"fb570",-- -1193
x"f71d0",-- -2275
x"f30c0",-- -3316
x"f0e40",-- -3868
x"f0f20",-- -3854
x"efe30",-- -4125
x"eca80",-- -4952
x"eaa80",-- -5464
x"ea470",-- -5561
x"ec560",-- -5034
x"ee7a0",-- -4486
x"f09b0",-- -3941
x"f2da0",-- -3366
x"f7b50",-- -2123
x"fe170",-- -489
x"024d0",-- 589
x"02c00",-- 704
x"02580",-- 600
x"032e0",-- 814
x"03e20",-- 994
x"02dc0",-- 732
x"ff790",-- -135
x"fc7d0",-- -899
x"fb3b0",-- -1221
x"fa550",-- -1451
x"f7e00",-- -2080
x"f5880",-- -2680
x"f5d30",-- -2605
x"f73e0",-- -2242
x"fa140",-- -1516
x"fddb0",-- -549
x"01670",-- 359
x"04730",-- 1139
x"073b0",-- 1851
x"09e20",-- 2530
x"0aae0",-- 2734
x"0ac20",-- 2754
x"0ab10",-- 2737
x"09fe0",-- 2558
x"09940",-- 2452
x"08340",-- 2100
x"05f80",-- 1528
x"02940",-- 660
x"ff560",-- -170
x"fd0e0",-- -754
x"fb1f0",-- -1249
x"f9ae0",-- -1618
x"f8e80",-- -1816
x"f8800",-- -1920
x"f9f40",-- -1548
x"fb590",-- -1191
x"fbec0",-- -1044
x"fbf80",-- -1032
x"fc350",-- -971
x"fe0a0",-- -502
x"fea20",-- -350
x"fead0",-- -339
x"ff510",-- -175
x"fff60",-- -10
x"013f0",-- 319
x"01a90",-- 425
x"01590",-- 345
x"00af0",-- 175
x"ff8a0",-- -118
x"ff800",-- -128
x"ff150",-- -235
x"ff470",-- -185
x"ffe20",-- -30
x"00c50",-- 197
x"02530",-- 595
x"04020",-- 1026
x"05920",-- 1426
x"063a0",-- 1594
x"07540",-- 1876
x"086d0",-- 2157
x"0a590",-- 2649
x"0c8e0",-- 3214
x"0f710",-- 3953
x"11ec0",-- 4588
x"12230",-- 4643
x"12610",-- 4705
x"11220",-- 4386
x"13400",-- 4928
x"16400",-- 5696
x"1b7d0",-- 7037
x"1ecc0",-- 7884
x"209a0",-- 8346
x"1f5b0",-- 8027
x"1c040",-- 7172
x"16910",-- 5777
x"0fb20",-- 4018
x"08580",-- 2136
x"fc410",-- -959
x"f5740",-- -2700
x"ef860",-- -4218
x"efba0",-- -4166
x"ee410",-- -4543
x"ed1b0",-- -4837
x"ec5a0",-- -5030
x"ef4c0",-- -4276
x"f3590",-- -3239
x"f4aa0",-- -2902
x"f7ea0",-- -2070
x"faaa0",-- -1366
x"fecb0",-- -309
x"ffc90",-- -55
x"011f0",-- 287
x"00700",-- 112
x"000d0",-- 13
x"fe7f0",-- -385
x"fd270",-- -729
x"fbf80",-- -1032
x"f92a0",-- -1750
x"f74d0",-- -2227
x"f51a0",-- -2790
x"f37a0",-- -3206
x"f1200",-- -3808
x"eef70",-- -4361
x"ec1c0",-- -5092
x"eae80",-- -5400
x"ec080",-- -5112
x"ec850",-- -4987
x"ee2b0",-- -4565
x"f1010",-- -3839
x"f4a50",-- -2907
x"f9950",-- -1643
x"fd6c0",-- -660
x"005c0",-- 92
x"013d0",-- 317
x"026b0",-- 619
x"033a0",-- 826
x"040f0",-- 1039
x"01e40",-- 484
x"fe6c0",-- -404
x"fd270",-- -729
x"fc080",-- -1016
x"fb020",-- -1278
x"f8050",-- -2043
x"f5e90",-- -2583
x"f6980",-- -2408
x"f9770",-- -1673
x"fc320",-- -974
x"fecb0",-- -309
x"01a60",-- 422
x"04db0",-- 1243
x"08770",-- 2167
x"0a930",-- 2707
x"0ae30",-- 2787
x"091a0",-- 2330
x"08ed0",-- 2285
x"08f00",-- 2288
x"08d40",-- 2260
x"07b50",-- 1973
x"04280",-- 1064
x"02f20",-- 754
x"01da0",-- 474
x"ff010",-- -255
x"faa20",-- -1374
x"f7e40",-- -2076
x"f8030",-- -2045
x"f9ab0",-- -1621
x"fadf0",-- -1313
x"fbbd0",-- -1091
x"fccd0",-- -819
x"fda40",-- -604
x"feaa0",-- -342
x"fe620",-- -414
x"fd100",-- -752
x"fbf60",-- -1034
x"fc7f0",-- -897
x"feda0",-- -294
x"00b20",-- 178
x"01a60",-- 422
x"01210",-- 289
x"01360",-- 310
x"01310",-- 305
x"00170",-- 23
x"fea00",-- -352
x"fda30",-- -605
x"fecf0",-- -305
x"00890",-- 137
x"020f0",-- 527
x"02be0",-- 702
x"03040",-- 772
x"03130",-- 787
x"031c0",-- 796
x"036a0",-- 874
x"03b20",-- 946
x"05860",-- 1414
x"08c00",-- 2240
x"0e5e0",-- 3678
x"12c20",-- 4802
x"15dd0",-- 5597
x"16550",-- 5717
x"13470",-- 4935
x"13720",-- 4978
x"12c50",-- 4805
x"16de0",-- 5854
x"1a810",-- 6785
x"1dad0",-- 7597
x"1f230",-- 7971
x"1f5b0",-- 8027
x"1c780",-- 7288
x"15af0",-- 5551
x"0d9c0",-- 3484
x"00440",-- 68
x"f47d0",-- -2947
x"ea170",-- -5609
x"eae60",-- -5402
x"eb520",-- -5294
x"ec290",-- -5079
x"ee7f0",-- -4481
x"f39d0",-- -3171
x"f9160",-- -1770
x"fa4d0",-- -1459
x"f8b60",-- -1866
x"f74a0",-- -2230
x"fa320",-- -1486
x"fc870",-- -889
x"ff740",-- -140
x"012e0",-- 302
x"04070",-- 1031
x"03f80",-- 1016
x"02840",-- 644
x"ff8f0",-- -113
x"f9da0",-- -1574
x"f3c20",-- -3134
x"f0140",-- -4076
x"efb30",-- -4173
x"efa70",-- -4185
x"efa70",-- -4185
x"ef390",-- -4295
x"efa60",-- -4186
x"efdb0",-- -4133
x"ef330",-- -4301
x"ed720",-- -4750
x"edde0",-- -4642
x"f1560",-- -3754
x"f6c30",-- -2365
x"fc490",-- -951
x"015e0",-- 350
x"052e0",-- 1326
x"06020",-- 1538
x"05ba0",-- 1466
x"03330",-- 819
x"ffee0",-- -18
x"fb8d0",-- -1139
x"f89b0",-- -1893
x"f8890",-- -1911
x"f9d30",-- -1581
x"faeb0",-- -1301
x"fa3e0",-- -1474
x"fb6a0",-- -1174
x"fc1b0",-- -997
x"fd530",-- -685
x"fdc10",-- -575
x"ff440",-- -188
x"02620",-- 610
x"054a0",-- 1354
x"09680",-- 2408
x"0bc60",-- 3014
x"0d080",-- 3336
x"0af70",-- 2807
x"094c0",-- 2380
x"07b30",-- 1971
x"04e50",-- 1253
x"01e90",-- 489
x"ffd60",-- -42
x"ffbc0",-- -68
x"00120",-- 18
x"ffee0",-- -18
x"fd990",-- -615
x"fc910",-- -879
x"fb360",-- -1226
x"fa760",-- -1418
x"f98d0",-- -1651
x"f99c0",-- -1636
x"fb540",-- -1196
x"fc8f0",-- -881
x"fe9b0",-- -357
x"ff0e0",-- -242
x"ff270",-- -217
x"fe3e0",-- -450
x"fddb0",-- -549
x"fda30",-- -605
x"fd530",-- -685
x"fd4c0",-- -692
x"fe070",-- -505
x"ffe70",-- -25
x"01040",-- 260
x"01710",-- 369
x"004e0",-- 78
x"ffc90",-- -55
x"ff3b0",-- -197
x"fe500",-- -432
x"fdc90",-- -567
x"fdae0",-- -594
x"fe530",-- -429
x"ff940",-- -108
x"017c0",-- 380
x"03360",-- 822
x"048c0",-- 1164
x"06160",-- 1558
x"087d0",-- 2173
x"0ae10",-- 2785
x"0d590",-- 3417
x"0fab0",-- 4011
x"12910",-- 4753
x"14bd0",-- 5309
x"15790",-- 5497
x"14b60",-- 5302
x"15e90",-- 5609
x"18000",-- 6144
x"19510",-- 6481
x"1ad40",-- 6868
x"1ac50",-- 6853
x"1c360",-- 7222
x"17830",-- 6019
x"14de0",-- 5342
x"0f950",-- 3989
x"062a0",-- 1578
x"f9e00",-- -1568
x"ee5a0",-- -4518
x"eda10",-- -4703
x"ea870",-- -5497
x"eac30",-- -5437
x"eae40",-- -5404
x"f1b80",-- -3656
x"f9720",-- -1678
x"fce30",-- -797
x"fcfc0",-- -772
x"fc410",-- -959
x"fe000",-- -512
x"fc160",-- -1002
x"fd2a0",-- -726
x"fcf00",-- -784
x"fee80",-- -280
x"ffb20",-- -78
x"01350",-- 309
x"01e50",-- 485
x"fdb30",-- -589
x"f9130",-- -1773
x"f3f30",-- -3085
x"f2930",-- -3437
x"ef7c0",-- -4228
x"ed380",-- -4808
x"ec690",-- -5015
x"eda70",-- -4697
x"f0c00",-- -3904
x"f1f40",-- -3596
x"f2100",-- -3568
x"f27a0",-- -3462
x"f51f0",-- -2785
x"f74d0",-- -2227
x"f9940",-- -1644
x"fcad0",-- -851
x"ffc10",-- -63
x"02ed0",-- 749
x"04300",-- 1072
x"04320",-- 1074
x"01900",-- 400
x"ff350",-- -203
x"fc7f0",-- -897
x"f9e70",-- -1561
x"f8fd0",-- -1795
x"f8b60",-- -1866
x"fafd0",-- -1283
x"fc6e0",-- -914
x"ff450",-- -187
x"01450",-- 325
x"02d20",-- 722
x"02870",-- 647
x"03680",-- 872
x"04c00",-- 1216
x"05180",-- 1304
x"05d10",-- 1489
x"061b0",-- 1563
x"07f60",-- 2038
x"08fe0",-- 2302
x"089b0",-- 2203
x"067f0",-- 1663
x"053d0",-- 1341
x"03540",-- 852
x"00f50",-- 245
x"ff490",-- -183
x"fdb00",-- -592
x"fcff0",-- -769
x"fd1b0",-- -741
x"fd470",-- -697
x"fce60",-- -794
x"fcaa0",-- -854
x"fcb90",-- -839
x"fc0c0",-- -1012
x"fb900",-- -1136
x"fbb50",-- -1099
x"fb090",-- -1271
x"fb850",-- -1147
x"fc9d0",-- -867
x"fe0a0",-- -502
x"fe4e0",-- -434
x"fe140",-- -492
x"feeb0",-- -277
x"ff6d0",-- -147
x"ff540",-- -172
x"fef30",-- -269
x"feed0",-- -275
x"ff260",-- -218
x"ffe50",-- -27
x"00080",-- 8
x"fff40",-- -12
x"ff6d0",-- -147
x"fef20",-- -270
x"fe5d0",-- -419
x"fe190",-- -487
x"fda30",-- -605
x"fd220",-- -734
x"fe4d0",-- -435
x"00660",-- 102
x"02700",-- 624
x"04c30",-- 1219
x"07040",-- 1796
x"0a140",-- 2580
x"0d740",-- 3444
x"0fff0",-- 4095
x"11f60",-- 4598
x"14960",-- 5270
x"17710",-- 6001
x"17f50",-- 6133
x"16a90",-- 5801
x"16450",-- 5701
x"18460",-- 6214
x"1a610",-- 6753
x"1a2c0",-- 6700
x"18a00",-- 6304
x"16020",-- 5634
x"13bc0",-- 5052
x"120e0",-- 4622
x"08200",-- 2080
x"fb9e0",-- -1122
x"f1560",-- -3754
x"ee380",-- -4552
x"ebe80",-- -5144
x"e8f80",-- -5896
x"ead50",-- -5419
x"f0320",-- -4046
x"f7330",-- -2253
x"fabc0",-- -1348
x"fecb0",-- -309
x"ff290",-- -215
x"fecd0",-- -307
x"fd4a0",-- -694
x"fe7d0",-- -387
x"000c0",-- 12
x"fe6c0",-- -404
x"fe340",-- -460
x"00e10",-- 225
x"03ea0",-- 1002
x"ff2c0",-- -212
x"fae80",-- -1304
x"f7a80",-- -2136
x"f49b0",-- -2917
x"f1110",-- -3823
x"ed5c0",-- -4772
x"ea380",-- -5576
x"ea650",-- -5531
x"ee4b0",-- -4533
x"f0190",-- -4071
x"f1c50",-- -3643
x"f3dd0",-- -3107
x"f6dc0",-- -2340
x"f98f0",-- -1649
x"fc550",-- -939
x"fde00",-- -544
x"fe850",-- -379
x"00390",-- 57
x"03130",-- 787
x"047a0",-- 1146
x"02980",-- 664
x"006c0",-- 108
x"00170",-- 23
x"ff4a0",-- -182
x"fccf0",-- -817
x"f9680",-- -1688
x"f82b0",-- -2005
x"fa0d0",-- -1523
x"fc840",-- -892
x"fdcc0",-- -564
x"ff5d0",-- -163
x"027b0",-- 635
x"04d40",-- 1236
x"06b60",-- 1718
x"07150",-- 1813
x"05c40",-- 1476
x"05440",-- 1348
x"060f0",-- 1551
x"06b30",-- 1715
x"062a0",-- 1578
x"05790",-- 1401
x"05950",-- 1429
x"06250",-- 1573
x"051a0",-- 1306
x"02960",-- 662
x"ff360",-- -202
x"fd490",-- -695
x"fce40",-- -796
x"fb6d0",-- -1171
x"fa070",-- -1529
x"f9ba0",-- -1606
x"fb200",-- -1248
x"fc660",-- -922
x"fca50",-- -859
x"fbee0",-- -1042
x"fb070",-- -1273
x"fb5c0",-- -1188
x"fc120",-- -1006
x"fbf30",-- -1037
x"fbfd0",-- -1027
x"fcd70",-- -809
x"fee10",-- -287
x"00b20",-- 178
x"015e0",-- 350
x"00a80",-- 168
x"fff40",-- -12
x"ff6a0",-- -150
x"feb70",-- -329
x"fd160",-- -746
x"fb9e0",-- -1122
x"fb740",-- -1164
x"fc0f0",-- -1009
x"fca70",-- -857
x"fc7b0",-- -901
x"fc800",-- -896
x"fd420",-- -702
x"fe6b0",-- -405
x"ffa60",-- -90
x"00390",-- 57
x"01710",-- 369
x"03ce0",-- 974
x"069b0",-- 1691
x"09170",-- 2327
x"0ab40",-- 2740
x"0c950",-- 3221
x"0f510",-- 3921
x"11d70",-- 4567
x"13010",-- 4865
x"14230",-- 5155
x"15820",-- 5506
x"15b90",-- 5561
x"15e20",-- 5602
x"16140",-- 5652
x"17420",-- 5954
x"18360",-- 6198
x"18a20",-- 6306
x"17ad0",-- 6061
x"15530",-- 5459
x"11d50",-- 4565
x"0bb30",-- 2995
x"02a80",-- 680
x"f7db0",-- -2085
x"f0210",-- -4063
x"eb590",-- -5287
x"e9110",-- -5871
x"e8150",-- -6123
x"eab60",-- -5450
x"f1db0",-- -3621
x"fa6e0",-- -1426
x"ff290",-- -215
x"00b10",-- 177
x"02410",-- 577
x"02e10",-- 737
x"02070",-- 519
x"ff2b0",-- -213
x"fc440",-- -956
x"fc960",-- -874
x"ff630",-- -157
x"ffc60",-- -58
x"ff580",-- -168
x"fef20",-- -270
x"fcf70",-- -777
x"f97c0",-- -1668
x"f5450",-- -2747
x"efbd0",-- -4163
x"eaf20",-- -5390
x"e9150",-- -5867
x"e99d0",-- -5731
x"ebe80",-- -5144
x"eecd0",-- -4403
x"f28e0",-- -3442
x"f7d60",-- -2090
x"fc8c0",-- -884
x"fea20",-- -350
x"ff790",-- -135
x"ffee0",-- -18
x"00af0",-- 175
x"018a0",-- 394
x"01420",-- 322
x"018a0",-- 394
x"02440",-- 580
x"02b40",-- 692
x"02640",-- 612
x"012c0",-- 300
x"feff0",-- -257
x"fc9b0",-- -869
x"fb420",-- -1214
x"f99e0",-- -1634
x"fa070",-- -1529
x"f8ca0",-- -1846
x"fa3c0",-- -1476
x"fda10",-- -607
x"02280",-- 552
x"05bf0",-- 1471
x"07530",-- 1875
x"0a000",-- 2560
x"0b630",-- 2915
x"0d310",-- 3377
x"0a190",-- 2585
x"08ca0",-- 2250
x"065d0",-- 1629
x"058b0",-- 1419
x"01120",-- 274
x"ff110",-- -239
x"feac0",-- -340
x"fd270",-- -729
x"fd100",-- -752
x"f8d00",-- -1840
x"fa4b0",-- -1461
x"f9a60",-- -1626
x"f9bf0",-- -1601
x"f7da0",-- -2086
x"f7ee0",-- -2066
x"fa9e0",-- -1378
x"faaa0",-- -1366
x"fb9a0",-- -1126
x"fcb10",-- -847
x"febb0",-- -325
x"ff290",-- -215
x"ffce0",-- -50
x"ff880",-- -120
x"ff880",-- -120
x"ff630",-- -157
x"ff020",-- -254
x"fede0",-- -290
x"fdcb0",-- -565
x"fd8b0",-- -629
x"fc820",-- -894
x"fbb70",-- -1097
x"faed0",-- -1299
x"f9330",-- -1741
x"f8940",-- -1900
x"f82a0",-- -2006
x"f8ee0",-- -1810
x"f9a90",-- -1623
x"fa670",-- -1433
x"fd100",-- -752
x"fef70",-- -265
x"015b0",-- 347
x"02c00",-- 704
x"04190",-- 1049
x"05d50",-- 1493
x"077c0",-- 1916
x"08870",-- 2183
x"092c0",-- 2348
x"0a450",-- 2629
x"0b580",-- 2904
x"0bf40",-- 3060
x"0c020",-- 3074
x"0c9a0",-- 3226
x"0ca40",-- 3236
x"0ddd0",-- 3549
x"0eed0",-- 3821
x"102a0",-- 4138
x"10720",-- 4210
x"12340",-- 4660
x"14e50",-- 5349
x"17120",-- 5906
x"183b0",-- 6203
x"19a30",-- 6563
x"1ba10",-- 7073
x"19760",-- 6518
x"14500",-- 5200
x"0b830",-- 2947
x"01090",-- 265
x"f5b50",-- -2635
x"eb840",-- -5244
x"e5200",-- -6880
x"e2d00",-- -7472
x"e4cb0",-- -6965
x"ea380",-- -5576
x"f3970",-- -3177
x"fdee0",-- -530
x"03880",-- 904
x"05e20",-- 1506
x"07060",-- 1798
x"060f0",-- 1551
x"02340",-- 564
x"fd010",-- -767
x"fa050",-- -1531
x"fa570",-- -1449
x"fcd70",-- -809
x"fd8a0",-- -630
x"fe890",-- -375
x"fff80",-- -8
x"00570",-- 87
x"fd150",-- -747
x"f7ab0",-- -2133
x"f2640",-- -3484
x"edd60",-- -4650
x"ea5b0",-- -5541
x"e8190",-- -6119
x"e95b0",-- -5797
x"ebf90",-- -5127
x"f0d70",-- -3881
x"f6b60",-- -2378
x"fc260",-- -986
x"008c0",-- 140
x"033a0",-- 826
x"04c20",-- 1218
x"05590",-- 1369
x"05600",-- 1376
x"034c0",-- 844
x"02280",-- 552
x"02230",-- 547
x"02160",-- 534
x"01030",-- 259
x"000f0",-- 15
x"ff300",-- -208
x"fe320",-- -462
x"fc9e0",-- -866
x"fa3c0",-- -1476
x"f9770",-- -1673
x"f9920",-- -1646
x"faff0",-- -1281
x"fce90",-- -791
x"007a0",-- 122
x"04300",-- 1072
x"088c0",-- 2188
x"0afa0",-- 2810
x"0d4c0",-- 3404
x"0bc70",-- 3015
x"08af0",-- 2223
x"071f0",-- 1823
x"04e50",-- 1253
x"02750",-- 629
x"fdb50",-- -587
x"fd290",-- -727
x"fdd30",-- -557
x"fead0",-- -339
x"fcf30",-- -781
x"f9ec0",-- -1556
x"f8b10",-- -1871
x"f9c10",-- -1599
x"f7ec0",-- -2068
x"f6670",-- -2457
x"f5790",-- -2695
x"f86e0",-- -1938
x"fcad0",-- -851
x"fe0d0",-- -499
x"ff800",-- -128
x"ffc90",-- -55
x"03180",-- 792
x"028f0",-- 655
x"ffa60",-- -90
x"fd3a0",-- -710
x"fc260",-- -986
x"fb900",-- -1136
x"fa660",-- -1434
x"f9ec0",-- -1556
x"f9c60",-- -1594
x"faf20",-- -1294
x"fc430",-- -957
x"fd2f0",-- -721
x"fc0f0",-- -1009
x"fbc20",-- -1086
x"fc2d0",-- -979
x"fc8e0",-- -882
x"fbd60",-- -1066
x"fac80",-- -1336
x"fb8d0",-- -1139
x"fd6c0",-- -660
x"fee40",-- -284
x"ffa30",-- -93
x"003a0",-- 58
x"03010",-- 769
x"05880",-- 1416
x"06af0",-- 1711
x"06fa0",-- 1786
x"07c40",-- 1988
x"08a40",-- 2212
x"09030",-- 2307
x"08350",-- 2101
x"07ae0",-- 1966
x"08890",-- 2185
x"09fb0",-- 2555
x"0b1d0",-- 2845
x"0bc10",-- 3009
x"0d950",-- 3477
x"102c0",-- 4140
x"114c0",-- 4428
x"134c0",-- 4940
x"142c0",-- 5164
x"156c0",-- 5484
x"16a70",-- 5799
x"17e60",-- 6118
x"19940",-- 6548
x"19560",-- 6486
x"191c0",-- 6428
x"13310",-- 4913
x"07c70",-- 1991
x"fc1c0",-- -996
x"f25c0",-- -3492
x"ea320",-- -5582
x"e0170",-- -8169
x"dc230",-- -9181
x"e1930",-- -7789
x"eccf0",-- -4913
x"f68c0",-- -2420
x"fdb80",-- -584
x"070e0",-- 1806
x"0f380",-- 3896
x"10750",-- 4213
x"09a90",-- 2473
x"03990",-- 921
x"ff490",-- -183
x"fb270",-- -1241
x"f6d00",-- -2352
x"f6020",-- -2558
x"f8ee0",-- -1810
x"fd7e0",-- -642
x"01d30",-- 467
x"03760",-- 886
x"03510",-- 849
x"00a70",-- 167
x"fb6f0",-- -1169
x"f3cc0",-- -3124
x"ec730",-- -5005
x"e67e0",-- -6530
x"e3090",-- -7415
x"e3b60",-- -7242
x"e8df0",-- -5921
x"f0820",-- -3966
x"f8b60",-- -1866
x"01e50",-- 485
x"0a5f0",-- 2655
x"0fb20",-- 4018
x"10730",-- 4211
x"0dee0",-- 3566
x"0ab30",-- 2739
x"06230",-- 1571
x"009e0",-- 158
x"fb620",-- -1182
x"f9720",-- -1678
x"f9f40",-- -1548
x"fa7f0",-- -1409
x"fb680",-- -1176
x"fd7c0",-- -644
x"ffb80",-- -72
x"001c0",-- 28
x"ff860",-- -122
x"fec60",-- -314
x"fe730",-- -397
x"fe140",-- -492
x"fee40",-- -284
x"00a70",-- 167
x"037c0",-- 892
x"06af0",-- 1711
x"09710",-- 2417
x"0bf60",-- 3062
x"0c7d0",-- 3197
x"0b720",-- 2930
x"08910",-- 2193
x"05710",-- 1393
x"014c0",-- 332
x"fc5f0",-- -929
x"f8b90",-- -1863
x"f6cd0",-- -2355
x"f6080",-- -2552
x"f51f0",-- -2785
x"f7330",-- -2253
x"f9a30",-- -1629
x"fba10",-- -1119
x"fc1e0",-- -994
x"fdae0",-- -594
x"fe490",-- -439
x"faa70",-- -1369
x"fa6b0",-- -1429
x"f9330",-- -1741
x"fb250",-- -1243
x"f9ba0",-- -1606
x"fac00",-- -1344
x"fef30",-- -269
x"02640",-- 612
x"03e90",-- 1001
x"00fc0",-- 252
x"02af0",-- 687
x"018b0",-- 395
x"fd920",-- -622
x"f8ca0",-- -1846
x"f6fc0",-- -2308
x"f6a20",-- -2398
x"f6370",-- -2505
x"f6580",-- -2472
x"f7fb0",-- -2053
x"fadf0",-- -1313
x"fd2f0",-- -721
x"feaa0",-- -342
x"fede0",-- -290
x"ff970",-- -105
x"ffce0",-- -50
x"ff580",-- -168
x"ff440",-- -188
x"001e0",-- 30
x"01940",-- 404
x"036f0",-- 879
x"051a0",-- 1306
x"07f90",-- 2041
x"090d0",-- 2317
x"09bf0",-- 2495
x"096d0",-- 2413
x"087f0",-- 2175
x"07bd0",-- 1981
x"05600",-- 1376
x"040d0",-- 1037
x"04370",-- 1079
x"05900",-- 1424
x"06b40",-- 1716
x"08a90",-- 2217
x"0b8a0",-- 2954
x"0f270",-- 3879
x"10230",-- 4131
x"11cd0",-- 4557
x"12270",-- 4647
x"12c20",-- 4802
x"11f60",-- 4598
x"10c80",-- 4296
x"11300",-- 4400
x"11d00",-- 4560
x"138d0",-- 5005
x"16980",-- 5784
x"155f0",-- 5471
x"07c40",-- 1988
x"fe390",-- -455
x"f9680",-- -1688
x"f2b60",-- -3402
x"e3970",-- -7273
x"db7a0",-- -9350
x"e0a00",-- -8032
x"ecad0",-- -4947
x"f4550",-- -2987
x"f3c20",-- -3134
x"00b20",-- 178
x"10be0",-- 4286
x"13360",-- 4918
x"0a9a0",-- 2714
x"07900",-- 1936
x"07b00",-- 1968
x"047f0",-- 1151
x"fc8e0",-- -882
x"f5840",-- -2684
x"f84e0",-- -1970
x"fcda0",-- -806
x"fe260",-- -474
x"fcd70",-- -809
x"fe250",-- -475
x"ffad0",-- -83
x"fe350",-- -459
x"f7060",-- -2298
x"ef510",-- -4271
x"ebef0",-- -5137
x"e8640",-- -6044
x"e6500",-- -6576
x"e92a0",-- -5846
x"ee380",-- -4552
x"f6c00",-- -2368
x"01030",-- 259
x"0a450",-- 2629
x"11dc0",-- 4572
x"15b50",-- 5557
x"14de0",-- 5342
x"12960",-- 4758
x"0e040",-- 3588
x"03bf0",-- 959
x"fa2a0",-- -1494
x"f5220",-- -2782
x"f2f20",-- -3342
x"f0480",-- -4024
x"efa70",-- -4185
x"f4250",-- -3035
x"fc170",-- -1001
x"00cf0",-- 207
x"02300",-- 560
x"053d0",-- 1341
x"08000",-- 2048
x"07f10",-- 2033
x"04a20",-- 1186
x"01c70",-- 455
x"01cb0",-- 459
x"02c10",-- 705
x"02430",-- 579
x"02910",-- 657
x"05580",-- 1368
x"07b20",-- 1970
x"07d80",-- 2008
x"06ea0",-- 1770
x"053a0",-- 1338
x"01b20",-- 434
x"fde70",-- -537
x"f9db0",-- -1573
x"f6bb0",-- -2373
x"f41c0",-- -3044
x"f3840",-- -3196
x"f5a40",-- -2652
x"f86c0",-- -1940
x"fb480",-- -1208
x"fc710",-- -911
x"fdb50",-- -587
x"00050",-- 5
x"ffb50",-- -75
x"fdc70",-- -569
x"fb570",-- -1193
x"fba80",-- -1112
x"fcb40",-- -844
x"fc430",-- -957
x"fc430",-- -957
x"fd380",-- -712
x"002a0",-- 42
x"00af0",-- 175
x"fee40",-- -284
x"fd850",-- -635
x"fd1a0",-- -742
x"fc2f0",-- -977
x"f96a0",-- -1686
x"f71a0",-- -2278
x"f75c0",-- -2212
x"f8260",-- -2010
x"f8ca0",-- -1846
x"f9a90",-- -1623
x"fb800",-- -1152
x"fe3e0",-- -450
x"005a0",-- 90
x"014e0",-- 334
x"01cc0",-- 460
x"022b0",-- 555
x"029e0",-- 670
x"023a0",-- 570
x"01cc0",-- 460
x"01bd0",-- 445
x"02620",-- 610
x"03940",-- 916
x"04a90",-- 1193
x"05a10",-- 1441
x"06b10",-- 1713
x"07c90",-- 1993
x"08680",-- 2152
x"08260",-- 2086
x"07510",-- 1873
x"06e10",-- 1761
x"06f40",-- 1780
x"07720",-- 1906
x"076d0",-- 1901
x"07f40",-- 2036
x"097b0",-- 2427
x"0c430",-- 3139
x"0e200",-- 3616
x"0e980",-- 3736
x"0fbd0",-- 4029
x"10900",-- 4240
x"11710",-- 4465
x"0ff50",-- 4085
x"0f8f0",-- 3983
x"0f920",-- 3986
x"11360",-- 4406
x"0dda0",-- 3546
x"059a0",-- 1434
x"00a30",-- 163
x"fc3f0",-- -961
x"f6d20",-- -2350
x"ecc60",-- -4922
x"e9950",-- -5739
x"ea800",-- -5504
x"efd40",-- -4140
x"f2670",-- -3481
x"f4b60",-- -2890
x"fdb70",-- -585
x"05ab0",-- 1451
x"096c0",-- 2412
x"073d0",-- 1853
x"08200",-- 2080
x"07ba0",-- 1978
x"060a0",-- 1546
x"008a0",-- 138
x"fbf90",-- -1031
x"fb250",-- -1243
x"fa960",-- -1386
x"f9c70",-- -1593
x"f7fd0",-- -2051
x"f9400",-- -1728
x"fad70",-- -1321
x"fbda0",-- -1062
x"f9130",-- -1773
x"f7510",-- -2223
x"f6710",-- -2447
x"f4980",-- -2920
x"f2be0",-- -3394
x"f1bb0",-- -3653
x"f2d20",-- -3374
x"f5b00",-- -2640
x"fa050",-- -1531
x"fde40",-- -540
x"02ed0",-- 749
x"074e0",-- 1870
x"0a210",-- 2593
x"0ba10",-- 2977
x"0ad60",-- 2774
x"07cc0",-- 1996
x"040a0",-- 1034
x"00410",-- 65
x"fc2a0",-- -982
x"f85a0",-- -1958
x"f5e40",-- -2588
x"f6120",-- -2542
x"f80c0",-- -2036
x"f9bc0",-- -1604
x"fc250",-- -987
x"fff60",-- -10
x"03940",-- 916
x"05720",-- 1394
x"05cb0",-- 1483
x"05a80",-- 1448
x"059f0",-- 1439
x"04c00",-- 1216
x"02800",-- 640
x"00d20",-- 210
x"00c10",-- 193
x"00fc0",-- 252
x"00e40",-- 228
x"00a20",-- 162
x"016d0",-- 365
x"021e0",-- 542
x"01c10",-- 449
x"00660",-- 102
x"fee60",-- -282
x"fdb70",-- -585
x"fc190",-- -999
x"fa9d0",-- -1379
x"f8eb0",-- -1813
x"f8bb0",-- -1861
x"f93e0",-- -1730
x"fa250",-- -1499
x"fb7b0",-- -1157
x"fcdc0",-- -804
x"fe910",-- -367
x"fe980",-- -360
x"00260",-- 38
x"fdec0",-- -532
x"fd070",-- -761
x"fbf80",-- -1032
x"fb090",-- -1271
x"fa8a0",-- -1398
x"f8a30",-- -1885
x"fb130",-- -1261
x"fadc0",-- -1316
x"fda10",-- -607
x"fd250",-- -731
x"fd720",-- -654
x"ff5d0",-- -163
x"fe660",-- -410
x"fd950",-- -619
x"fb940",-- -1132
x"fb850",-- -1147
x"faf00",-- -1296
x"fa550",-- -1451
x"f9f10",-- -1551
x"fb070",-- -1273
x"fc9d0",-- -867
x"fe9b0",-- -357
x"fffe0",-- -2
x"019e0",-- 414
x"03ab0",-- 939
x"04940",-- 1172
x"05670",-- 1383
x"045f0",-- 1119
x"04530",-- 1107
x"03ec0",-- 1004
x"03040",-- 772
x"029b0",-- 667
x"023a0",-- 570
x"03120",-- 786
x"04430",-- 1091
x"05150",-- 1301
x"06730",-- 1651
x"08000",-- 2048
x"09ce0",-- 2510
x"0a7f0",-- 2687
x"0b490",-- 2889
x"0b7c0",-- 2940
x"0bb20",-- 2994
x"0b860",-- 2950
x"0b090",-- 2825
x"0ae00",-- 2784
x"0a110",-- 2577
x"0b220",-- 2850
x"0bc90",-- 3017
x"0d710",-- 3441
x"0ea50",-- 3749
x"10810",-- 4225
x"13ad0",-- 5037
x"0fd30",-- 4051
x"0a520",-- 2642
x"05fe0",-- 1534
x"01630",-- 355
x"f9f40",-- -1548
x"efb80",-- -4168
x"ecd90",-- -4903
x"ebf70",-- -5129
x"eeb70",-- -4425
x"ee980",-- -4456
x"f16b0",-- -3733
x"fb4a0",-- -1206
x"02570",-- 599
x"05800",-- 1408
x"06440",-- 1604
x"0abe0",-- 2750
x"0b900",-- 2960
x"09810",-- 2433
x"03fb0",-- 1019
x"00020",-- 2
x"fe7f0",-- -385
x"fb990",-- -1127
x"f80a0",-- -2038
x"f55c0",-- -2724
x"f7ae0",-- -2130
x"f9650",-- -1691
x"fa8a0",-- -1398
x"f9540",-- -1708
x"fad20",-- -1326
x"fc580",-- -936
x"fae40",-- -1308
x"f8190",-- -2023
x"f6280",-- -2520
x"f6530",-- -2477
x"f6070",-- -2553
x"f5df0",-- -2593
x"f6660",-- -2458
x"fab40",-- -1356
x"feff0",-- -257
x"01d80",-- 472
x"04db0",-- 1243
x"080f0",-- 2063
x"09e00",-- 2528
x"091c0",-- 2332
x"07630",-- 1891
x"04980",-- 1176
x"018b0",-- 395
x"fd9a0",-- -614
x"f9f30",-- -1549
x"f81c0",-- -2020
x"f6f80",-- -2312
x"f7150",-- -2283
x"f8710",-- -1935
x"fb680",-- -1176
x"fe700",-- -400
x"01810",-- 385
x"03e40",-- 996
x"06500",-- 1616
x"07a60",-- 1958
x"06ea0",-- 1770
x"05bd0",-- 1469
x"04990",-- 1177
x"03330",-- 819
x"00c00",-- 192
x"ff300",-- -208
x"fe940",-- -364
x"fee60",-- -282
x"fed40",-- -300
x"fec50",-- -315
x"ffdf0",-- -33
x"00da0",-- 218
x"00cb0",-- 203
x"ffb50",-- -75
x"fed40",-- -300
x"fde00",-- -544
x"fc690",-- -919
x"fa5c0",-- -1444
x"f91f0",-- -1761
x"f93e0",-- -1730
x"f9d60",-- -1578
x"fa9e0",-- -1378
x"fc7f0",-- -897
x"ff020",-- -254
x"019c0",-- 412
x"03a40",-- 932
x"04d60",-- 1238
x"05530",-- 1363
x"05170",-- 1303
x"037e0",-- 894
x"006b0",-- 107
x"fd9c0",-- -612
x"fa750",-- -1419
x"f8070",-- -2041
x"f5ba0",-- -2630
x"f4bc0",-- -2884
x"f5090",-- -2807
x"f6710",-- -2447
x"f8530",-- -1965
x"f9e20",-- -1566
x"fc940",-- -876
x"fe5a0",-- -422
x"ffd30",-- -45
x"005d0",-- 93
x"00930",-- 147
x"00ac0",-- 172
x"002f0",-- 47
x"ffb80",-- -72
x"ff580",-- -168
x"ffe50",-- -27
x"fffe0",-- -2
x"00960",-- 150
x"01290",-- 297
x"01f90",-- 505
x"025f0",-- 607
x"022f0",-- 559
x"020d0",-- 525
x"014c0",-- 332
x"00a30",-- 163
x"ff590",-- -167
x"fea80",-- -344
x"fe6c0",-- -404
x"fe4e0",-- -434
x"fed40",-- -300
x"ffa90",-- -87
x"00f00",-- 240
x"026e0",-- 622
x"03920",-- 914
x"047b0",-- 1147
x"05920",-- 1426
x"059c0",-- 1436
x"05e00",-- 1504
x"05810",-- 1409
x"05e20",-- 1506
x"05e50",-- 1509
x"06250",-- 1573
x"07220",-- 1826
x"07900",-- 1936
x"09450",-- 2373
x"0a000",-- 2560
x"0b440",-- 2884
x"0ba80",-- 2984
x"0c7f0",-- 3199
x"0cd20",-- 3282
x"0cc00",-- 3264
x"0ca90",-- 3241
x"0c570",-- 3159
x"0c7a0",-- 3194
x"0b860",-- 2950
x"0b290",-- 2857
x"09620",-- 2402
x"06cd0",-- 1741
x"033d0",-- 829
x"00210",-- 33
x"fc8a0",-- -886
x"f8030",-- -2045
x"f5160",-- -2794
x"f32c0",-- -3284
x"f32e0",-- -3282
x"f3ae0",-- -3154
x"f4e60",-- -2842
x"f7ce0",-- -2098
x"fc8a0",-- -886
x"00280",-- 40
x"02820",-- 642
x"05510",-- 1361
x"07ec0",-- 2028
x"08d20",-- 2258
x"07e40",-- 2020
x"067d0",-- 1661
x"04a70",-- 1191
x"02d10",-- 721
x"ffcc0",-- -52
x"fc9d0",-- -867
x"fa6e0",-- -1426
x"f9330",-- -1741
x"f80a0",-- -2038
x"f6be0",-- -2370
x"f6390",-- -2503
x"f6c60",-- -2362
x"f7310",-- -2255
x"f71b0",-- -2277
x"f72f0",-- -2257
x"f7b00",-- -2128
x"f8760",-- -1930
x"f92a0",-- -1750
x"f9850",-- -1659
x"fa850",-- -1403
x"fc760",-- -906
x"fe3a0",-- -454
x"ff720",-- -142
x"00dc0",-- 220
x"02960",-- 662
x"036f0",-- 879
x"03760",-- 886
x"02d10",-- 721
x"01f90",-- 505
x"00ac0",-- 172
x"feb10",-- -335
x"fcca0",-- -822
x"fb420",-- -1214
x"fa4e0",-- -1458
x"f9bf0",-- -1601
x"fa110",-- -1519
x"fb1b0",-- -1253
x"fcd50",-- -811
x"fee10",-- -287
x"00e10",-- 225
x"031c0",-- 796
x"049e0",-- 1182
x"05760",-- 1398
x"05940",-- 1428
x"054c0",-- 1356
x"042a0",-- 1066
x"026b0",-- 619
x"00f00",-- 240
x"ff6d0",-- -147
x"fe5f0",-- -417
x"fd5e0",-- -674
x"fd060",-- -762
x"fd530",-- -685
x"fdf90",-- -519
x"fea30",-- -349
x"ff180",-- -232
x"ffe20",-- -30
x"00480",-- 72
x"00480",-- 72
x"ff9f0",-- -97
x"ff1a0",-- -230
x"feaa0",-- -342
x"fe0d0",-- -499
x"fd770",-- -649
x"fd670",-- -665
x"fdfd0",-- -515
x"feb20",-- -334
x"ff8f0",-- -113
x"00570",-- 87
x"01590",-- 345
x"02050",-- 517
x"02370",-- 567
x"01a90",-- 425
x"00f90",-- 249
x"ffee0",-- -18
x"fe980",-- -360
x"fce40",-- -796
x"fbb30",-- -1101
x"f8fa0",-- -1798
x"f8260",-- -2010
x"f8300",-- -2000
x"f77f0",-- -2177
x"f7920",-- -2158
x"f7b30",-- -2125
x"faeb0",-- -1301
x"fb880",-- -1144
x"fd220",-- -734
x"fddd0",-- -547
x"ff3b0",-- -197
x"01c20",-- 450
x"00ac0",-- 172
x"007d0",-- 125
x"009d0",-- 157
x"016f0",-- 367
x"00a30",-- 163
x"ff540",-- -172
x"ff270",-- -217
x"ff800",-- -128
x"ff4f0",-- -177
x"fed20",-- -302
x"fe660",-- -410
x"fefa0",-- -262
x"003c0",-- 60
x"fff90",-- -7
x"003f0",-- 63
x"007a0",-- 122
x"01c20",-- 450
x"02430",-- 579
x"01ab0",-- 427
x"02390",-- 569
x"030b0",-- 779
x"04620",-- 1122
x"04f90",-- 1273
x"05790",-- 1401
x"06ea0",-- 1770
x"08f40",-- 2292
x"0a080",-- 2568
x"0a400",-- 2624
x"0b4f0",-- 2895
x"0c820",-- 3202
x"0d680",-- 3432
x"0ceb0",-- 3307
x"0d0e0",-- 3342
x"0d6a0",-- 3434
x"0df30",-- 3571
x"0e130",-- 3603
x"0e2d0",-- 3629
x"0f630",-- 3939
x"105a0",-- 4186
x"103c0",-- 4156
x"0eae0",-- 3758
x"09830",-- 2435
x"03b70",-- 951
x"00980",-- 152
x"fa6c0",-- -1428
x"f2da0",-- -3366
x"ecff0",-- -4865
x"ed930",-- -4717
x"edf90",-- -4615
x"edd40",-- -4652
x"efbb0",-- -4165
x"f41e0",-- -3042
x"fd3a0",-- -710
x"01060",-- 262
x"02780",-- 632
x"05fb0",-- 1531
x"0c310",-- 3121
x"0cf50",-- 3317
x"09f80",-- 2552
x"08530",-- 2131
x"07860",-- 1926
x"069a0",-- 1690
x"01950",-- 405
x"fd1f0",-- -737
x"fb0c0",-- -1268
x"fb290",-- -1239
x"f8700",-- -1936
x"f4ed0",-- -2835
x"f3390",-- -3271
x"f3b00",-- -3152
x"f4300",-- -3024
x"f1a70",-- -3673
x"f0bc0",-- -3908
x"f2870",-- -3449
x"f4d20",-- -2862
x"f59a0",-- -2662
x"f6620",-- -2462
x"f8df0",-- -1825
x"fd760",-- -650
x"01210",-- 289
x"01cc0",-- 460
x"03b70",-- 951
x"07150",-- 1813
x"08cd0",-- 2253
x"07b50",-- 1973
x"05f30",-- 1523
x"05270",-- 1319
x"04200",-- 1056
x"01540",-- 340
x"fd2f0",-- -721
x"fb590",-- -1191
x"fa870",-- -1401
x"f9470",-- -1721
x"f7fe0",-- -2050
x"f8300",-- -2000
x"fa2f0",-- -1489
x"fc820",-- -894
x"fe2a0",-- -470
x"00070",-- 7
x"03470",-- 839
x"05900",-- 1424
x"069a0",-- 1690
x"073d0",-- 1853
x"07ae0",-- 1966
x"07420",-- 1858
x"060d0",-- 1549
x"047b0",-- 1147
x"02d90",-- 729
x"01380",-- 312
x"ff770",-- -137
x"fe3c0",-- -452
x"fd9c0",-- -612
x"fcda0",-- -806
x"fc4e0",-- -946
x"fc760",-- -906
x"fd1a0",-- -742
x"fd450",-- -699
x"fd2e0",-- -722
x"fd850",-- -635
x"fe370",-- -457
x"fe8c0",-- -372
x"fdf80",-- -520
x"fe690",-- -407
x"ff3b0",-- -197
x"ffe70",-- -25
x"00050",-- 5
x"00730",-- 115
x"01860",-- 390
x"02390",-- 569
x"02640",-- 612
x"01ad0",-- 429
x"01b00",-- 432
x"01470",-- 327
x"001e0",-- 30
x"fe780",-- -392
x"fd130",-- -749
x"fc2d0",-- -979
x"faff0",-- -1281
x"fa190",-- -1511
x"f9400",-- -1728
x"f9df0",-- -1569
x"fab20",-- -1358
x"fba10",-- -1119
x"fcc60",-- -826
x"fe580",-- -424
x"00840",-- 132
x"01fd0",-- 509
x"03530",-- 851
x"03ec0",-- 1004
x"050d0",-- 1293
x"05360",-- 1334
x"04d70",-- 1239
x"03f40",-- 1012
x"03170",-- 791
x"026c0",-- 620
x"013f0",-- 319
x"003f0",-- 63
x"ff3d0",-- -195
x"ff2e0",-- -210
x"fed40",-- -300
x"febc0",-- -324
x"feb60",-- -330
x"ff170",-- -233
x"ffb50",-- -75
x"ffd50",-- -43
x"ffd60",-- -42
x"ffdb0",-- -37
x"fff30",-- -13
x"ffce0",-- -50
x"ffa10",-- -95
x"ff8d0",-- -115
x"ffce0",-- -50
x"00340",-- 52
x"00bb0",-- 187
x"013f0",-- 319
x"01e20",-- 482
x"02980",-- 664
x"03090",-- 777
x"03440",-- 836
x"033f0",-- 831
x"02c60",-- 710
x"024d0",-- 589
x"018d0",-- 397
x"005a0",-- 90
x"ff240",-- -220
x"fe1b0",-- -485
x"fd810",-- -639
x"fce30",-- -797
x"fc9e0",-- -866
x"fce80",-- -792
x"fdbd0",-- -579
x"febe0",-- -322
x"ff710",-- -143
x"00440",-- 68
x"013f0",-- 319
x"01d50",-- 469
x"01c20",-- 450
x"01540",-- 340
x"00fc0",-- 252
x"009e0",-- 158
x"fff10",-- -15
x"ff310",-- -207
x"ff4c0",-- -180
x"ff800",-- -128
x"ffee0",-- -18
x"00870",-- 135
x"01650",-- 357
x"026b0",-- 619
x"031a0",-- 794
x"03a60",-- 934
x"03920",-- 914
x"03830",-- 899
x"02ea0",-- 746
x"01fd0",-- 509
x"00cf0",-- 207
x"ffc10",-- -63
x"fef30",-- -269
x"fe460",-- -442
x"fde40",-- -540
x"fde70",-- -537
x"fe7a0",-- -390
x"ff2b0",-- -213
x"00080",-- 8
x"00c80",-- 200
x"019f0",-- 415
x"02410",-- 577
x"027b0",-- 635
x"02480",-- 584
x"01ec0",-- 492
x"016d0",-- 365
x"00ac0",-- 172
x"ffc90",-- -55
x"ff040",-- -252
x"fe6b0",-- -405
x"fe210",-- -479
x"fe140",-- -492
x"fe430",-- -445
x"fe9e0",-- -354
x"ff360",-- -202
x"ffe20",-- -30
x"005f0",-- 95
x"00b60",-- 182
x"00e80",-- 232
x"01060",-- 262
x"00d40",-- 212
x"00840",-- 132
x"ffe70",-- -25
x"ff8b0",-- -117
x"ff1c0",-- -228
x"feaf0",-- -337
x"fe5a0",-- -422
x"fe4d0",-- -435
x"fe8c0",-- -372
x"feb40",-- -332
x"fefa0",-- -262
x"ff440",-- -188
x"ffd00",-- -48
x"001b0",-- 27
x"004d0",-- 77
x"00530",-- 83
x"00670",-- 103
x"00730",-- 115
x"003e0",-- 62
x"00000",-- 0
x"ffbc0",-- -68
x"ffb80",-- -72
x"ff880",-- -120
x"ff800",-- -128
x"ff720",-- -142
x"ff970",-- -105
x"ff100",-- -240
x"fefc0",-- -260
x"fef30",-- -269
x"fe7a0",-- -390
x"fdf40",-- -524
x"fd590",-- -679
x"fd8b0",-- -629
x"fcca0",-- -822
x"fc820",-- -894
x"fbf80",-- -1032
x"fbe20",-- -1054
x"fc640",-- -924
x"fc000",-- -1024
x"fc280",-- -984
x"fce60",-- -794
x"fdf90",-- -519
x"fe6e0",-- -402
x"fee10",-- -287
x"ffc60",-- -58
x"00980",-- 152
x"00eb0",-- 235
x"00e80",-- 232
x"00dc0",-- 220
x"00f50",-- 245
x"00eb0",-- 235
x"002a0",-- 42
x"ffb70",-- -73
x"ff470",-- -185
x"ff2e0",-- -210
x"fee80",-- -280
x"fe930",-- -365
x"fee80",-- -280
x"ff260",-- -218
x"ff950",-- -107
x"00070",-- 7
x"006b0",-- 107
x"00dc0",-- 220
x"01830",-- 387
x"01f90",-- 505
x"023e0",-- 574
x"02980",-- 664
x"03210",-- 801
x"038a0",-- 906
x"03c70",-- 967
x"04200",-- 1056
x"04750",-- 1141
x"05310",-- 1329
x"05670",-- 1383
x"05b30",-- 1459
x"06140",-- 1556
x"06700",-- 1648
x"06900",-- 1680
x"068b0",-- 1675
x"069f0",-- 1695
x"06a50",-- 1701
x"06ae0",-- 1710
x"067a0",-- 1658
x"06840",-- 1668
x"067a0",-- 1658
x"06410",-- 1601
x"057c0",-- 1404
x"04f90",-- 1273
x"03fb0",-- 1019
x"02980",-- 664
x"013d0",-- 317
x"ffd50",-- -43
x"fe990",-- -359
x"fd510",-- -687
x"fc5f0",-- -929
x"fbc60",-- -1082
x"fba10",-- -1119
x"fb9a0",-- -1126
x"fba80",-- -1112
x"fc410",-- -959
x"fd2e0",-- -722
x"fdc10",-- -575
x"fe3f0",-- -449
x"ff010",-- -255
x"ffbd0",-- -67
x"000c0",-- 12
x"00000",-- 0
x"000f0",-- 15
x"00080",-- 8
x"ffc90",-- -55
x"ff240",-- -220
x"fe960",-- -362
x"fe140",-- -492
x"fd670",-- -665
x"fc7f0",-- -897
x"fb9a0",-- -1126
x"fb090",-- -1271
x"fa710",-- -1423
x"f9bf0",-- -1601
x"f9570",-- -1705
x"f9540",-- -1708
x"f9940",-- -1644
x"f9df0",-- -1569
x"fa5c0",-- -1444
x"fb250",-- -1243
x"fc230",-- -989
x"fd150",-- -747
x"fe0d0",-- -499
x"ff060",-- -250
x"fff60",-- -10
x"00af0",-- 175
x"01100",-- 272
x"01590",-- 345
x"01600",-- 352
x"01710",-- 369
x"011f0",-- 287
x"00d90",-- 217
x"00800",-- 128
x"00250",-- 37
x"ffe50",-- -27
x"ff9c0",-- -100
x"ff720",-- -142
x"ff5d0",-- -163
x"ff7c0",-- -132
x"ff8d0",-- -115
x"ffb20",-- -78
x"ffe90",-- -23
x"00300",-- 48
x"00760",-- 118
x"00ad0",-- 173
x"00c50",-- 197
x"00fa0",-- 250
x"011a0",-- 282
x"01380",-- 312
x"01420",-- 322
x"01400",-- 320
x"014a0",-- 330
x"01380",-- 312
x"011a0",-- 282
x"00d90",-- 217
x"00b60",-- 182
x"00690",-- 105
x"000d0",-- 13
x"ffb50",-- -75
x"ff5d0",-- -163
x"ff010",-- -255
x"fecb0",-- -309
x"fea80",-- -344
x"fe840",-- -380
x"fe930",-- -365
x"fead0",-- -339
x"fee10",-- -287
x"ff110",-- -239
x"ff540",-- -172
x"ff920",-- -110
x"ffdb0",-- -37
x"00000",-- 0
x"fffd0",-- -3
x"ffe90",-- -23
x"ffe40",-- -28
x"ffc20",-- -62
x"ff880",-- -120
x"ff450",-- -187
x"ff150",-- -235
x"fef00",-- -272
x"febe0",-- -322
x"fe9e0",-- -354
x"fe930",-- -365
x"fead0",-- -339
x"fecb0",-- -309
x"feed0",-- -275
x"ff300",-- -208
x"ff800",-- -128
x"ffe50",-- -27
x"00370",-- 55
x"008c0",-- 140
x"00df0",-- 223
x"011f0",-- 287
x"01560",-- 342
x"016f0",-- 367
x"01860",-- 390
x"01800",-- 384
x"01580",-- 344
x"01270",-- 295
x"010d0",-- 269
x"00d00",-- 208
x"00a80",-- 168
x"007d0",-- 125
x"00660",-- 102
x"00530",-- 83
x"003a0",-- 58
x"00480",-- 72
x"00320",-- 50
x"003c0",-- 60
x"004e0",-- 78
x"004b0",-- 75
x"004b0",-- 75
x"00570",-- 87
x"00620",-- 98
x"00570",-- 87
x"00620",-- 98
x"005f0",-- 95
x"00610",-- 97
x"00660",-- 102
x"00750",-- 117
x"00850",-- 133
x"00990",-- 153
x"00a80",-- 168
x"00ac0",-- 172
x"00ca0",-- 202
x"00c50",-- 197
x"00c60",-- 198
x"00b70",-- 183
x"00ac0",-- 172
x"00870",-- 135
x"004e0",-- 78
x"002b0",-- 43
x"fffe0",-- -2
x"ffda0",-- -38
x"ffa30",-- -93
x"ff920",-- -110
x"ff900",-- -112
x"ff810",-- -127
x"ff7c0",-- -132
x"ff8d0",-- -115
x"ffad0",-- -83
x"ffd00",-- -48
x"00000",-- 0
x"00440",-- 68
x"00a70",-- 167
x"00ef0",-- 239
x"01270",-- 295
x"01670",-- 359
x"019a0",-- 410
x"01b00",-- 432
x"01ab0",-- 427
x"01ad0",-- 429
x"01a10",-- 417
x"01790",-- 377
x"01530",-- 339
x"01220",-- 290
x"00f00",-- 240
x"00b60",-- 182
x"00840",-- 132
x"005d0",-- 93
x"00440",-- 68
x"002a0",-- 42
x"00190",-- 25
x"00230",-- 35
x"00250",-- 37
x"002a0",-- 42
x"00370",-- 55
x"00460",-- 70
x"00640",-- 100
x"00710",-- 113
x"00800",-- 128
x"00870",-- 135
x"008c0",-- 140
x"00840",-- 132
x"00760",-- 118
x"00710",-- 113
x"004e0",-- 78
x"00320",-- 50
x"000c0",-- 12
x"fff10",-- -15
x"ffbf0",-- -65
x"ff950",-- -107
x"ff790",-- -135
x"ff5b0",-- -165
x"ff510",-- -175
x"ff3b0",-- -197
x"ff420",-- -190
x"ff3a0",-- -198
x"ff4e0",-- -178
x"ff510",-- -175
x"ff5b0",-- -165
x"ff6c0",-- -148
x"ff6d0",-- -147
x"ff810",-- -127
x"ff710",-- -143
x"ff6d0",-- -147
x"ff6c0",-- -148
x"ff670",-- -153
x"ff650",-- -155
x"ff680",-- -152
x"ff6f0",-- -145
x"ff790",-- -135
x"ff7c0",-- -132
x"ff8d0",-- -115
x"ff970",-- -105
x"ff920",-- -110
x"ff990",-- -103
x"ff950",-- -107
x"ff9c0",-- -100
x"ff8d0",-- -115
x"ff880",-- -120
x"ff810",-- -127
x"ff740",-- -140
x"ff710",-- -143
x"ff5d0",-- -163
x"ff580",-- -168
x"ff670",-- -153
x"ff6d0",-- -147
x"ff740",-- -140
x"ff880",-- -120
x"ff950",-- -107
x"ffa30",-- -93
x"ff100",-- -240
x"fef70",-- -265
x"fea50",-- -347
x"fe570",-- -425
x"fd9f0",-- -609
x"fd160",-- -746
x"fd530",-- -685
x"fd110",-- -751
x"fd470",-- -697
x"fd200",-- -736
x"fdfe0",-- -514
x"fecf0",-- -305
x"ff400",-- -192
x"ffb70",-- -73
x"00370",-- 55
x"013a0",-- 314
x"016c0",-- 364
x"016a0",-- 362
x"01580",-- 344
x"018a0",-- 394
x"01620",-- 354
x"00d20",-- 210
x"00370",-- 55
x"ffdb0",-- -37
x"ffb00",-- -80
x"ff1c0",-- -228
x"fea30",-- -349
x"fe5d0",-- -419
x"fe8a0",-- -374
x"fe9b0",-- -357
x"fe850",-- -379
x"fed70",-- -297
x"ff490",-- -183
x"ffd10",-- -47
x"002f0",-- 47
x"00960",-- 150
x"01240",-- 292
x"01ba0",-- 442
x"02280",-- 552
x"02500",-- 592
x"02870",-- 647
x"02bc0",-- 700
x"02d70",-- 727
x"02960",-- 662
x"02410",-- 577
x"02050",-- 517
x"01f30",-- 499
x"019f0",-- 415
x"01260",-- 294
x"00eb0",-- 235
x"00e80",-- 232
x"00e10",-- 225
x"00960",-- 150
x"00a00",-- 160
x"00d50",-- 213
x"01220",-- 290
x"011f0",-- 287
x"01360",-- 310
x"018a0",-- 394
x"01c40",-- 452
x"01ce0",-- 462
x"019f0",-- 415
x"01cc0",-- 460
x"01d00",-- 464
x"01b70",-- 439
x"01620",-- 354
x"012e0",-- 302
x"010b0",-- 267
x"00cb0",-- 203
x"00960",-- 150
x"00530",-- 83
x"006c0",-- 108
x"00550",-- 85
x"004b0",-- 75
x"004e0",-- 78
x"00690",-- 105
x"00730",-- 115
x"004e0",-- 78
x"00690",-- 105
x"005f0",-- 95
x"00530",-- 83
x"00260",-- 38
x"001b0",-- 27
x"002a0",-- 42
x"fff90",-- -7
x"ffdf0",-- -33
x"ffcb0",-- -53
x"ffd50",-- -43
x"ffda0",-- -38
x"ffb50",-- -75
x"ffa30",-- -93
x"ffad0",-- -83
x"ff9c0",-- -100
x"ff6d0",-- -147
x"ff540",-- -172
x"ff600",-- -160
x"ff4e0",-- -178
x"ff330",-- -205
x"ff220",-- -222
x"ff0c0",-- -244
x"ff210",-- -223
x"ff180",-- -232
x"ff0c0",-- -244
x"ff1f0",-- -225
x"ff2b0",-- -213
x"ff400",-- -192
x"ff380",-- -200
x"ff300",-- -208
x"ff330",-- -205
x"ff2e0",-- -210
x"ff180",-- -232
x"fef30",-- -269
x"fede0",-- -290
x"febb0",-- -325
x"fea20",-- -350
x"fe7a0",-- -390
x"fe570",-- -425
x"fe340",-- -460
x"fe3c0",-- -452
x"fe3e0",-- -450
x"fe3e0",-- -450
x"fe550",-- -427
x"fe5c0",-- -420
x"fe7d0",-- -387
x"fe7d0",-- -387
x"fe990",-- -359
x"fea20",-- -350
x"fea80",-- -344
x"feaa0",-- -342
x"fe9b0",-- -357
x"fea30",-- -349
x"fea50",-- -347
x"febc0",-- -324
x"feaf0",-- -337
x"feb70",-- -329
x"fed40",-- -300
x"fee80",-- -280
x"ff0c0",-- -244
x"ff220",-- -222
x"ff470",-- -185
x"ff6f0",-- -145
x"ff830",-- -125
x"ff970",-- -105
x"ffae0",-- -82
x"ffc60",-- -58
x"ffc60",-- -58
x"ffd50",-- -43
x"ffd60",-- -42
x"fff10",-- -15
x"ffee0",-- -18
x"000c0",-- 12
x"002a0",-- 42
x"00430",-- 67
x"00750",-- 117
x"00960",-- 150
x"00e10",-- 225
x"00e10",-- 225
x"011c0",-- 284
x"01380",-- 312
x"01710",-- 369
x"01a30",-- 419
x"01c90",-- 457
x"02260",-- 550
x"02490",-- 585
x"02b20",-- 690
x"03130",-- 787
x"03810",-- 897
x"04170",-- 1047
x"04870",-- 1159
x"05440",-- 1348
x"05d80",-- 1496
x"06900",-- 1680
x"071d0",-- 1821
x"07e40",-- 2020
x"08af0",-- 2223
x"08ca0",-- 2250
x"06a20",-- 1698
x"051a0",-- 1306
x"04490",-- 1097
x"01510",-- 337
x"fd4f0",-- -689
x"f9fe0",-- -1538
x"f9830",-- -1661
x"f70e0",-- -2290
x"f4e90",-- -2839
x"f3930",-- -3181
x"f4570",-- -2985
x"f6bb0",-- -2373
x"f6dc0",-- -2340
x"f7cb0",-- -2101
x"fa440",-- -1468
x"fe700",-- -400
x"fff60",-- -10
x"00ca0",-- 202
x"02d70",-- 727
x"053d0",-- 1341
x"06410",-- 1601
x"04ed0",-- 1261
x"04620",-- 1122
x"04160",-- 1046
x"03a10",-- 929
x"011d0",-- 285
x"fe620",-- -414
x"fccf0",-- -817
x"fbc10",-- -1087
x"f9da0",-- -1574
x"f75b0",-- -2213
x"f6cb0",-- -2357
x"f6c80",-- -2360
x"f6d00",-- -2352
x"f6d70",-- -2345
x"f7590",-- -2215
x"f8c30",-- -1853
x"fa9d0",-- -1379
x"fc550",-- -939
x"fd1a0",-- -742
x"febe0",-- -322
x"00b90",-- 185
x"020c0",-- 524
x"026e0",-- 622
x"02bc0",-- 700
x"036a0",-- 874
x"03e00",-- 992
x"03990",-- 921
x"02a30",-- 675
x"02710",-- 625
x"025c0",-- 604
x"020a0",-- 522
x"00fa0",-- 250
x"00500",-- 80
x"00850",-- 133
x"00610",-- 97
x"ffdf0",-- -33
x"ff530",-- -173
x"ffce0",-- -50
x"001b0",-- 27
x"fff90",-- -7
x"ffd50",-- -43
x"001b0",-- 27
x"00b60",-- 182
x"00cb0",-- 203
x"00c50",-- 197
x"00eb0",-- 235
x"016d0",-- 365
x"01990",-- 409
x"01710",-- 369
x"01900",-- 400
x"01bf0",-- 447
x"01cc0",-- 460
x"019a0",-- 410
x"01790",-- 377
x"014a0",-- 330
x"00fc0",-- 252
x"00960",-- 150
x"00480",-- 72
x"fff60",-- -10
x"ff5d0",-- -163
x"ff240",-- -220
x"fef20",-- -270
x"fedc0",-- -292
x"fea00",-- -352
x"feb20",-- -334
x"ff020",-- -254
x"ff4a0",-- -182
x"ff800",-- -128
x"ff790",-- -135
x"fffe0",-- -2
x"005a0",-- 90
x"006b0",-- 107
x"00440",-- 68
x"005c0",-- 92
x"00850",-- 133
x"00320",-- 50
x"ffbf0",-- -65
x"ff6a0",-- -150
x"ff650",-- -155
x"ff310",-- -207
x"fed50",-- -299
x"fe9e0",-- -354
x"feda0",-- -294
x"ff1c0",-- -228
x"ff180",-- -232
x"ff4c0",-- -180
x"ffbf0",-- -65
x"00640",-- 100
x"00a80",-- 168
x"00d90",-- 217
x"01380",-- 312
x"019a0",-- 410
x"01c90",-- 457
x"01bf0",-- 447
x"01ae0",-- 430
x"01a30",-- 419
x"019c0",-- 412
x"01450",-- 325
x"01030",-- 259
x"00d70",-- 215
x"00c00",-- 192
x"008e0",-- 142
x"00490",-- 73
x"000f0",-- 15
x"fff40",-- -12
x"ffe20",-- -30
x"ffb50",-- -75
x"ff900",-- -112
x"ff6d0",-- -147
x"ff770",-- -137
x"ff6c0",-- -148
x"ff740",-- -140
x"ff800",-- -128
x"ffae0",-- -82
x"fffb0",-- -5
x"002f0",-- 47
x"00530",-- 83
x"009b0",-- 155
x"00e90",-- 233
x"012b0",-- 299
x"014f0",-- 335
x"01450",-- 325
x"014c0",-- 332
x"01290",-- 297
x"01030",-- 259
x"00960",-- 150
x"004e0",-- 78
x"00000",-- 0
x"ffbf0",-- -65
x"ff6d0",-- -147
x"ff1c0",-- -228
x"ff100",-- -240
x"fefd0",-- -259
x"ff010",-- -255
x"fef00",-- -272
x"fefd0",-- -259
x"ff2b0",-- -213
x"ff620",-- -158
x"ff860",-- -122
x"ff9c0",-- -100
x"fff80",-- -8
x"00370",-- 55
x"00750",-- 117
x"00aa0",-- 170
x"01040",-- 260
x"01600",-- 352
x"01970",-- 407
x"01c70",-- 455
x"01db0",-- 475
x"02050",-- 517
x"01fe0",-- 510
x"01df0",-- 479
x"01990",-- 409
x"016c0",-- 364
x"012e0",-- 302
x"00c50",-- 197
x"00670",-- 103
x"00250",-- 37
x"00000",-- 0
x"ffc90",-- -55
x"ff990",-- -103
x"ff7c0",-- -132
x"ff8a0",-- -118
x"ffa30",-- -93
x"ffbc0",-- -68
x"ffcc0",-- -52
x"000f0",-- 15
x"00410",-- 65
x"00570",-- 87
x"006b0",-- 107
x"00840",-- 132
x"00980",-- 152
x"00850",-- 133
x"006b0",-- 107
x"004e0",-- 78
x"003c0",-- 60
x"00120",-- 18
x"fff80",-- -8
x"ffea0",-- -22
x"ffdb0",-- -37
x"ffd60",-- -42
x"ffce0",-- -50
x"ffd50",-- -43
x"ffc70",-- -57
x"ffbf0",-- -65
x"ffbd0",-- -67
x"ffbd0",-- -67
x"ffb70",-- -73
x"ff8f0",-- -113
x"ff760",-- -138
x"ff630",-- -157
x"ff4e0",-- -178
x"ff100",-- -240
x"ff070",-- -249
x"ff110",-- -239
x"ff270",-- -217
x"ff260",-- -218
x"ff3d0",-- -195
x"ff830",-- -125
x"ffa90",-- -87
x"ffdd0",-- -35
x"fff90",-- -7
x"003f0",-- 63
x"00640",-- 100
x"006b0",-- 107
x"00640",-- 100
x"005c0",-- 92
x"005d0",-- 93
x"002f0",-- 47
x"fffe0",-- -2
x"ffc20",-- -62
x"ffb20",-- -78
x"ff800",-- -128
x"ff580",-- -168
x"ff420",-- -190
x"ff4a0",-- -182
x"ff590",-- -167
x"ff580",-- -168
x"ff7b0",-- -133
x"ff8a0",-- -118
x"ffb20",-- -78
x"ffc90",-- -55
x"ffe70",-- -25
x"fff80",-- -8
x"fff60",-- -10
x"000a0",-- 10
x"00000",-- 0
x"fff90",-- -7
x"ffe50",-- -27
x"ffd10",-- -47
x"ffc60",-- -58
x"ffb80",-- -72
x"ffa30",-- -93
x"ff9f0",-- -97
x"ffab0",-- -85
x"ffa90",-- -87
x"ffb20",-- -78
x"ffab0",-- -85
x"ffc60",-- -58
x"ffcb0",-- -53
x"ffcc0",-- -52
x"ffc60",-- -58
x"ffc20",-- -62
x"ffbc0",-- -68
x"ffa10",-- -95
x"ff830",-- -125
x"ff710",-- -143
x"ff670",-- -153
x"ff580",-- -168
x"ff580",-- -168
x"ff580",-- -168
x"ff830",-- -125
x"ff990",-- -103
x"ffc60",-- -58
x"ffee0",-- -18
x"00200",-- 32
x"00670",-- 103
x"007a0",-- 122
x"00a30",-- 163
x"00ac0",-- 172
x"00b60",-- 182
x"00a80",-- 168
x"00730",-- 115
x"00430",-- 67
x"00170",-- 23
x"fff10",-- -15
x"ffad0",-- -83
x"ff7c0",-- -132
x"ff600",-- -160
x"ff4f0",-- -177
x"ff400",-- -192
x"ff4e0",-- -178
x"ff710",-- -143
x"ffb20",-- -78
x"ffe20",-- -30
x"00070",-- 7
x"004e0",-- 78
x"00870",-- 135
x"00b20",-- 178
x"00bb0",-- 187
x"00bc0",-- 188
x"00b90",-- 185
x"00a70",-- 167
x"00870",-- 135
x"00480",-- 72
x"000a0",-- 10
x"ffe70",-- -25
x"ffa90",-- -87
x"ff850",-- -123
x"ff600",-- -160
x"ff600",-- -160
x"ff760",-- -138
x"ff790",-- -135
x"ff860",-- -122
x"ffad0",-- -83
x"ffe50",-- -27
x"00050",-- 5
x"00280",-- 40
x"00460",-- 70
x"004b0",-- 75
x"003e0",-- 62
x"00340",-- 52
x"000c0",-- 12
x"fff10",-- -15
x"ffd80",-- -40
x"ffbc0",-- -68
x"ff9c0",-- -100
x"ff830",-- -125
x"ff790",-- -135
x"ff800",-- -128
x"ff900",-- -112
x"ff9c0",-- -100
x"ffb70",-- -73
x"ffe40",-- -28
x"00000",-- 0
x"00030",-- 3
x"000f0",-- 15
x"00230",-- 35
x"003f0",-- 63
x"00250",-- 37
x"00190",-- 25
x"00020",-- 2
x"fff40",-- -12
x"fff80",-- -8
x"ffea0",-- -22
x"ffdb0",-- -37
x"ffdb0",-- -37
x"fff80",-- -8
x"ffee0",-- -18
x"fff40",-- -12
x"ffb00",-- -80
x"ffab0",-- -85
x"ffa90",-- -87
x"ff470",-- -185
x"fef70",-- -265
x"fe6c0",-- -404
x"fe7f0",-- -385
x"fe0f0",-- -497
x"fdae0",-- -594
x"fd880",-- -632
x"fd560",-- -682
x"fdc20",-- -574
x"fd760",-- -650
x"fd8b0",-- -629
x"fdd80",-- -552
x"fe1e0",-- -482
x"fe800",-- -384
x"fe710",-- -399
x"fef50",-- -267
x"ff5d0",-- -163
x"ffb20",-- -78
x"ffd30",-- -45
x"ffe90",-- -23
x"003a0",-- 58
x"00490",-- 73
x"003a0",-- 58
x"00160",-- 22
x"00080",-- 8
x"00000",-- 0
x"ffe00",-- -32
x"ff9f0",-- -97
x"ffa40",-- -92
x"ffa60",-- -90
x"ffb20",-- -78
x"ffce0",-- -50
x"ffe20",-- -30
x"002f0",-- 47
x"00780",-- 120
x"00eb0",-- 235
x"01220",-- 290
x"01770",-- 375
x"01e90",-- 489
x"02390",-- 569
x"027b0",-- 635
x"028e0",-- 654
x"02c60",-- 710
x"03010",-- 769
x"03010",-- 769
x"03010",-- 769
x"03040",-- 772
x"03450",-- 837
x"036d0",-- 877
x"03740",-- 884
x"03900",-- 912
x"03b80",-- 952
x"040a0",-- 1034
x"041b0",-- 1051
x"042d0",-- 1069
x"045f0",-- 1119
x"048e0",-- 1166
x"04be0",-- 1214
x"04910",-- 1169
x"049e0",-- 1182
x"04940",-- 1172
x"04750",-- 1141
x"03fb0",-- 1019
x"037e0",-- 894
x"03040",-- 772
x"023c0",-- 572
x"01720",-- 370
x"008f0",-- 143
x"ffd50",-- -43
x"ff040",-- -252
x"fe340",-- -460
x"fd9e0",-- -610
x"fd1b0",-- -741
x"fccf0",-- -817
x"fc7f0",-- -897
x"fc7a0",-- -902
x"fc930",-- -877
x"fcd40",-- -812
x"fd1d0",-- -739
x"fd720",-- -654
x"fe050",-- -507
x"fe5c0",-- -420
x"fec10",-- -319
x"fed20",-- -302
x"ff010",-- -255
x"ff100",-- -240
x"fecf0",-- -305
x"fe7a0",-- -390
x"fe190",-- -487
x"fdc90",-- -567
x"fd340",-- -716
x"fcb20",-- -846
x"fc3f0",-- -961
x"fbef0",-- -1041
x"fba80",-- -1112
x"fb6c0",-- -1172
x"fb670",-- -1177
x"fb810",-- -1151
x"fbd10",-- -1071
x"fc210",-- -991
x"fc910",-- -879
x"fd0c0",-- -756
x"fd900",-- -624
x"fe110",-- -495
x"fe760",-- -394
x"fed90",-- -295
x"ff310",-- -207
x"ff920",-- -110
x"ffce0",-- -50
x"ffee0",-- -18
x"00000",-- 0
x"000c0",-- 12
x"00230",-- 35
x"00140",-- 20
x"001b0",-- 27
x"00280",-- 40
x"003a0",-- 58
x"00460",-- 70
x"00530",-- 83
x"00760",-- 118
x"008f0",-- 143
x"00ac0",-- 172
x"00be0",-- 190
x"00c00",-- 192
x"00d70",-- 215
x"00e90",-- 233
x"00d20",-- 210
x"00c80",-- 200
x"00be0",-- 190
x"00b40",-- 180
x"008e0",-- 142
x"00760",-- 118
x"00640",-- 100
x"00530",-- 83
x"00550",-- 85
x"00320",-- 50
x"001b0",-- 27
x"000f0",-- 15
x"00250",-- 37
x"001b0",-- 27
x"00110",-- 17
x"000f0",-- 15
x"00020",-- 2
x"fffe0",-- -2
x"ffef0",-- -17
x"ffee0",-- -18
x"ffce0",-- -50
x"ffc60",-- -58
x"ffa80",-- -88
x"ff810",-- -127
x"ff6f0",-- -145
x"ff760",-- -138
x"ff670",-- -153
x"ff400",-- -192
x"ff4a0",-- -182
x"ff470",-- -185
x"ff3a0",-- -198
x"ff350",-- -203
x"ff350",-- -203
x"ff3d0",-- -195
x"ff4e0",-- -178
x"ff4e0",-- -178
x"ff4e0",-- -178
x"ff6a0",-- -150
x"ff830",-- -125
x"ffa60",-- -90
x"ffa90",-- -87
x"ffc20",-- -62
x"ffe20",-- -30
x"fff10",-- -15
x"00190",-- 25
x"00160",-- 22
x"003e0",-- 62
x"00570",-- 87
x"00690",-- 105
x"00840",-- 132
x"007d0",-- 125
x"009d0",-- 157
x"00940",-- 148
x"009b0",-- 155
x"00a20",-- 162
x"009d0",-- 157
x"00a30",-- 163
x"007f0",-- 127
x"00840",-- 132
x"00730",-- 115
x"00730",-- 115
x"00690",-- 105
x"004d0",-- 77
x"003f0",-- 63
x"00390",-- 57
x"00440",-- 68
x"00260",-- 38
x"002d0",-- 45
x"00230",-- 35
x"002a0",-- 42
x"00250",-- 37
x"00210",-- 33
x"002d0",-- 45
x"00300",-- 48
x"00410",-- 65
x"005a0",-- 90
x"00640",-- 100
x"00620",-- 98
x"00750",-- 117
x"00700",-- 112
x"00760",-- 118
x"005d0",-- 93
x"004e0",-- 78
x"00410",-- 65
x"002b0",-- 43
x"00170",-- 23
x"fffd0",-- -3
x"fff60",-- -10
x"ffec0",-- -20
x"ffe20",-- -30
x"ffd60",-- -42
x"ffdb0",-- -37
x"ffe90",-- -23
x"fff60",-- -10
x"00000",-- 0
x"00120",-- 18
x"002b0",-- 43
x"00440",-- 68
x"00320",-- 50
x"002b0",-- 43
x"00280",-- 40
x"00080",-- 8
x"00000",-- 0
x"ffe40",-- -28
x"ffdf0",-- -33
x"ffc40",-- -60
x"ffb70",-- -73
x"ffbc0",-- -68
x"ff9f0",-- -97
x"ffc10",-- -63
x"ffc10",-- -63
x"ffbd0",-- -67
x"ffd00",-- -48
x"ffc60",-- -58
x"ffdf0",-- -33
x"ffd10",-- -47
x"ffdb0",-- -37
x"ffce0",-- -50
x"ffb80",-- -72
x"ffb20",-- -78
x"ff8d0",-- -115
x"ff800",-- -128
x"ff670",-- -153
x"ff350",-- -203
x"ff1d0",-- -227
x"ff0c0",-- -244
x"ff070",-- -249
x"fef20",-- -270
x"ff040",-- -252
x"ff150",-- -235
x"ff1d0",-- -227
x"ff3b0",-- -197
x"ff530",-- -173
x"ff920",-- -110
x"ffb50",-- -75
x"ffd50",-- -43
x"000c0",-- 12
x"002f0",-- 47
x"00580",-- 88
x"00640",-- 100
x"00850",-- 133
x"00a30",-- 163
x"00a50",-- 165
x"00a30",-- 163
x"00980",-- 152
x"00a30",-- 163
x"00990",-- 153
x"00730",-- 115
x"00710",-- 113
x"006b0",-- 107
x"006c0",-- 108
x"00520",-- 82
x"00520",-- 82
x"00700",-- 112
x"008a0",-- 138
x"009e0",-- 158
x"00ac0",-- 172
x"00d20",-- 210
x"00ef0",-- 239
x"010d0",-- 269
x"012b0",-- 299
x"01360",-- 310
x"014c0",-- 332
x"01420",-- 322
x"01510",-- 337
x"01360",-- 310
x"01180",-- 280
x"00f70",-- 247
x"00df0",-- 223
x"00da0",-- 218
x"00a20",-- 162
x"00890",-- 137
x"007b0",-- 123
x"006e0",-- 110
x"005d0",-- 93
x"002a0",-- 42
x"00280",-- 40
x"001b0",-- 27
x"00210",-- 33
x"00120",-- 18
x"00000",-- 0
x"00080",-- 8
x"fff80",-- -8
x"fff80",-- -8
x"ffd50",-- -43
x"ffbd0",-- -67
x"ffb30",-- -77
x"ffa60",-- -90
x"ff8a0",-- -118
x"ff710",-- -143
x"ff5b0",-- -165
x"ff5d0",-- -163
x"ff400",-- -192
x"ff240",-- -220
x"ff0e0",-- -242
x"ff020",-- -254
x"ff0b0",-- -245
x"fefa0",-- -262
x"fef50",-- -267
x"ff010",-- -255
x"ff060",-- -250
x"ff020",-- -254
x"ff040",-- -252
x"fefc0",-- -260
x"fefd0",-- -259
x"ff010",-- -255
x"fef50",-- -267
x"fef30",-- -269
x"ff060",-- -250
x"ff1d0",-- -227
x"ff1c0",-- -228
x"ff300",-- -208
x"ff470",-- -185
x"ff5d0",-- -163
x"ff760",-- -138
x"ff770",-- -137
x"ff900",-- -112
x"ffa30",-- -93
x"ffb80",-- -72
x"ffc90",-- -55
x"ffd50",-- -43
x"ffd80",-- -40
x"ffd80",-- -40
x"ffd30",-- -45
x"ffdf0",-- -33
x"ffe50",-- -27
x"ffec0",-- -20
x"fff10",-- -15
x"ffe90",-- -23
x"ffee0",-- -18
x"fff30",-- -13
x"fff80",-- -8
x"00000",-- 0
x"001c0",-- 28
x"00340",-- 52
x"004d0",-- 77
x"00690",-- 105
x"00800",-- 128
x"00a30",-- 163
x"00bc0",-- 188
x"00d40",-- 212
x"00d70",-- 215
x"00c30",-- 195
x"00bc0",-- 188
x"00a80",-- 168
x"00930",-- 147
x"007d0",-- 125
x"007a0",-- 122
x"006c0",-- 108
x"005a0",-- 90
x"005a0",-- 90
x"00530",-- 83
x"00550",-- 85
x"00620",-- 98
x"00730",-- 115
x"008e0",-- 142
x"00990",-- 153
x"00b90",-- 185
x"00bc0",-- 188
x"00c00",-- 192
x"00bc0",-- 188
x"00a50",-- 165
x"00820",-- 130
x"00670",-- 103
x"00570",-- 87
x"00350",-- 53
x"00370",-- 55
x"00350",-- 53
x"002b0",-- 43
x"00320",-- 50
x"00530",-- 83
x"00670",-- 103
x"00690",-- 105
x"00660",-- 102
x"00710",-- 113
x"006b0",-- 107
x"00530",-- 83
x"002b0",-- 43
x"000c0",-- 12
x"001e0",-- 30
x"fff10",-- -15
x"fff80",-- -8
x"ffea0",-- -22
x"fffe0",-- -2
x"ffe50",-- -27
x"ffdd0",-- -35
x"00030",-- 3
x"fffd0",-- -3
x"ffe70",-- -25
x"ffc20",-- -62
x"ffce0",-- -50
x"ffbc0",-- -68
x"ff6d0",-- -147
x"ff400",-- -192
x"ff130",-- -237
x"ff100",-- -240
x"feb90",-- -327
x"fe730",-- -397
x"fe520",-- -430
x"fe700",-- -400
x"fe730",-- -397
x"fe440",-- -444
x"fe5c0",-- -420
x"fe760",-- -394
x"feac0",-- -340
x"fe8c0",-- -372
x"fe730",-- -397
x"feb70",-- -329
x"feb20",-- -334
x"feaf0",-- -337
x"fe890",-- -375
x"feaa0",-- -342
x"feda0",-- -294
x"febe0",-- -322
x"fea80",-- -344
x"feb90",-- -327
x"feeb0",-- -277
x"fede0",-- -290
x"fed00",-- -304
x"fef70",-- -265
x"ff180",-- -232
x"ff2b0",-- -213
x"ff380",-- -200
x"ff4a0",-- -182
x"ff830",-- -125
x"ffa60",-- -90
x"ffd10",-- -47
x"ffe00",-- -32
x"00080",-- 8
x"003e0",-- 62
x"006b0",-- 107
x"008f0",-- 143
x"00af0",-- 175
x"00d40",-- 212
x"00f70",-- 247
x"012c0",-- 300
x"012b0",-- 299
x"011f0",-- 287
x"01470",-- 327
x"015b0",-- 347
x"01420",-- 322
x"01360",-- 310
x"015d0",-- 349
x"018a0",-- 394
x"019a0",-- 410
x"01a10",-- 417
x"01d00",-- 464
x"020d0",-- 525
x"02210",-- 545
x"02350",-- 565
x"023e0",-- 574
x"02320",-- 562
x"025f0",-- 607
x"02750",-- 629
x"026c0",-- 620
x"02850",-- 645
x"02bc0",-- 700
x"02be0",-- 702
x"02980",-- 664
x"027f0",-- 639
x"028c0",-- 652
x"02940",-- 660
x"02750",-- 629
x"022b0",-- 555
x"02230",-- 547
x"02530",-- 595
x"023c0",-- 572
x"02480",-- 584
x"024b0",-- 587
x"026b0",-- 619
x"02690",-- 617
x"02390",-- 569
x"022f0",-- 559
x"02050",-- 517
x"02070",-- 519
x"01ba0",-- 442
x"01860",-- 390
x"01530",-- 339
x"01290",-- 297
x"014c0",-- 332
x"01100",-- 272
x"00c50",-- 197
x"00840",-- 132
x"008c0",-- 140
x"00370",-- 55
x"ff710",-- -143
x"ff1c0",-- -228
x"fec00",-- -320
x"fe820",-- -382
x"fe020",-- -510
x"fda10",-- -607
x"fd8d0",-- -627
x"fd8a0",-- -630
x"fda40",-- -604
x"fd3d0",-- -707
x"fd4f0",-- -689
x"fd760",-- -650
x"fd8d0",-- -627
x"fd650",-- -667
x"fd360",-- -714
x"fd470",-- -697
x"fd4f0",-- -689
x"fd420",-- -702
x"fcbc0",-- -836
x"fc7b0",-- -901
x"fc980",-- -872
x"fc6c0",-- -916
x"fc340",-- -972
x"fc110",-- -1007
x"fc670",-- -921
x"fca70",-- -857
x"fcb40",-- -844
x"fccb0",-- -821
x"fcf00",-- -784
x"fd3a0",-- -710
x"fd360",-- -714
x"fd200",-- -736
x"fd1a0",-- -742
x"fd330",-- -717
x"fd580",-- -680
x"fd270",-- -729
x"fd200",-- -736
x"fd4c0",-- -692
x"fd9c0",-- -612
x"fdcc0",-- -564
x"fde20",-- -542
x"fe170",-- -489
x"fe5c0",-- -420
x"fea50",-- -347
x"fea20",-- -350
x"fea50",-- -347
x"fee80",-- -280
x"ff1a0",-- -230
x"ff350",-- -203
x"ff3b0",-- -197
x"ff590",-- -167
x"ffb20",-- -78
x"ffe50",-- -27
x"00000",-- 0
x"00250",-- 37
x"00850",-- 133
x"00cf0",-- 207
x"00e40",-- 228
x"01100",-- 272
x"011a0",-- 282
x"011f0",-- 287
x"010b0",-- 267
x"00f70",-- 247
x"00e40",-- 228
x"00c00",-- 192
x"00c00",-- 192
x"00bc0",-- 188
x"00bb0",-- 187
x"00fa0",-- 250
x"012b0",-- 299
x"01650",-- 357
x"018d0",-- 397
x"01d50",-- 469
x"02080",-- 520
x"02210",-- 545
x"02580",-- 600
x"02760",-- 630
x"02670",-- 615
x"024b0",-- 587
x"02670",-- 615
x"02870",-- 647
x"026b0",-- 619
x"024b0",-- 587
x"02500",-- 592
x"02490",-- 585
x"023c0",-- 572
x"024b0",-- 587
x"02430",-- 579
x"02440",-- 580
x"024d0",-- 589
x"02570",-- 599
x"02620",-- 610
x"02550",-- 597
x"02690",-- 617
x"02800",-- 640
x"02760",-- 630
x"024b0",-- 587
x"02430",-- 579
x"02780",-- 632
x"02a20",-- 674
x"02be0",-- 702
x"029b0",-- 667
x"02910",-- 657
x"02a70",-- 679
x"02780",-- 632
x"02080",-- 520
x"01bf0",-- 447
x"01530",-- 339
x"00d40",-- 212
x"00490",-- 73
x"ffd10",-- -47
x"ff7c0",-- -132
x"ff290",-- -215
x"fefa0",-- -262
x"fe800",-- -384
x"fe5a0",-- -422
x"fe3a0",-- -454
x"fe2d0",-- -467
x"fe200",-- -480
x"fdce0",-- -562
x"fe0a0",-- -502
x"fe0c0",-- -500
x"fdfd0",-- -515
x"fe030",-- -509
x"fe1c0",-- -484
x"fe4b0",-- -437
x"fe4e0",-- -434
x"fe530",-- -429
x"fe190",-- -487
x"fe030",-- -509
x"fda80",-- -600
x"fd3a0",-- -710
x"fce90",-- -791
x"fc820",-- -894
x"fc820",-- -894
x"fc490",-- -951
x"fc3f0",-- -961
x"fc710",-- -911
x"fcc50",-- -827
x"fd1d0",-- -739
x"fd530",-- -685
x"fdc40",-- -572
x"fdfd0",-- -515
x"fe620",-- -414
x"fe890",-- -375
x"fe9b0",-- -357
x"fec50",-- -315
x"fed90",-- -295
x"fef80",-- -264
x"fee40",-- -284
x"ff070",-- -249
x"ff1f0",-- -225
x"ff3f0",-- -193
x"ff790",-- -135
x"ff830",-- -125
x"ff9e0",-- -98
x"ffa30",-- -93
x"ffad0",-- -83
x"ffb80",-- -72
x"ffcc0",-- -52
x"ffee0",-- -18
x"fff80",-- -8
x"00120",-- 18
x"003f0",-- 63
x"00760",-- 118
x"00990",-- 153
x"00d50",-- 213
x"011a0",-- 282
x"01260",-- 294
x"013f0",-- 319
x"016c0",-- 364
x"018d0",-- 397
x"017e0",-- 382
x"01830",-- 387
x"01720",-- 370
x"011f0",-- 287
x"00e90",-- 233
x"00bb0",-- 187
x"009b0",-- 155
x"00730",-- 115
x"00670",-- 103
x"005f0",-- 95
x"00750",-- 117
x"007b0",-- 123
x"00940",-- 148
x"009d0",-- 157
x"006b0",-- 107
x"004b0",-- 75
x"00390",-- 57
x"00280",-- 40
x"000c0",-- 12
x"ffe50",-- -27
x"ffe50",-- -27
x"ffdf0",-- -33
x"ffbc0",-- -68
x"ffae0",-- -82
x"ffba0",-- -70
x"ffc20",-- -62
x"ffc90",-- -55
x"ffdd0",-- -35
x"00050",-- 5
x"00170",-- 23
x"00430",-- 67
x"00990",-- 153
x"00b40",-- 180
x"00cf0",-- 207
x"00bc0",-- 188
x"00a20",-- 162
x"00660",-- 102
x"00280",-- 40
x"000d0",-- 13
x"ffd10",-- -47
x"ffc60",-- -58
x"ffda0",-- -38
x"ffe20",-- -30
x"ff9c0",-- -100
x"ff880",-- -120
x"ffb00",-- -80
x"ffa40",-- -92
x"ffba0",-- -70
x"ffba0",-- -70
x"ffd80",-- -40
x"fffd0",-- -3
x"00250",-- 37
x"003f0",-- 63
x"00610",-- 97
x"00ad0",-- 173
x"00cb0",-- 203
x"00a00",-- 160
x"00670",-- 103
x"005d0",-- 93
x"005d0",-- 93
x"00080",-- 8
x"ffce0",-- -50
x"ffc20",-- -62
x"ff990",-- -103
x"ff740",-- -140
x"ff6a0",-- -150
x"ff600",-- -160
x"ff740",-- -140
x"ff900",-- -112
x"ff530",-- -173
x"ff240",-- -220
x"ff6d0",-- -147
x"ff940",-- -108
x"ff920",-- -110
x"ff850",-- -123
x"ffa40",-- -92
x"fff30",-- -13
x"fffd0",-- -3
x"ffdb0",-- -37
x"ffe20",-- -30
x"000a0",-- 10
x"00140",-- 20
x"ffd50",-- -43
x"ffa60",-- -90
x"ffad0",-- -83
x"ff860",-- -122
x"ff4e0",-- -178
x"ff330",-- -205
x"ff2b0",-- -213
x"ff180",-- -232
x"ff240",-- -220
x"ff4a0",-- -182
x"ff510",-- -175
x"ff790",-- -135
x"ffbf0",-- -65
x"ffee0",-- -18
x"00020",-- 2
x"fffe0",-- -2
x"00390",-- 57
x"00480",-- 72
x"00210",-- 33
x"00140",-- 20
x"00200",-- 32
x"00490",-- 73
x"00350",-- 53
x"00530",-- 83
x"00700",-- 112
x"00a00",-- 160
x"00cf0",-- 207
x"00c00",-- 192
x"00e30",-- 227
x"00e80",-- 232
x"00e40",-- 228
x"00de0",-- 222
x"00e30",-- 227
x"00fc0",-- 252
x"00e40",-- 228
x"00e60",-- 230
x"00f20",-- 242
x"00eb0",-- 235
x"00eb0",-- 235
x"00c00",-- 192
x"00cb0",-- 203
x"01100",-- 272
x"01060",-- 262
x"00cb0",-- 203
x"00eb0",-- 235
x"01560",-- 342
x"013b0",-- 315
x"00e80",-- 232
x"00eb0",-- 235
x"01220",-- 290
x"00fa0",-- 250
x"00930",-- 147
x"00820",-- 130
x"007a0",-- 122
x"004b0",-- 75
x"004e0",-- 78
x"00490",-- 73
x"00480",-- 72
x"007d0",-- 125
x"00a50",-- 165
x"007d0",-- 125
x"00700",-- 112
x"00a00",-- 160
x"00be0",-- 190
x"00960",-- 150
x"00440",-- 68
x"00170",-- 23
x"00170",-- 23
x"00050",-- 5
x"ffc20",-- -62
x"ff770",-- -137
x"ff770",-- -137
x"ff850",-- -123
x"ff5d0",-- -163
x"ff150",-- -235
x"ff0e0",-- -242
x"ff2e0",-- -210
x"ff090",-- -247
x"feda0",-- -294
x"fec10",-- -319
x"fec10",-- -319
x"fef20",-- -270
x"fefa0",-- -262
x"fef30",-- -269
x"ff220",-- -222
x"ff5d0",-- -163
x"ff710",-- -143
x"ff6d0",-- -147
x"ff790",-- -135
x"ff7b0",-- -133
x"ff860",-- -122
x"ff9c0",-- -100
x"ffa80",-- -88
x"ffce0",-- -50
x"000d0",-- 13
x"00430",-- 67
x"00460",-- 70
x"00570",-- 87
x"00690",-- 105
x"00520",-- 82
x"00030",-- 3
x"ffa60",-- -90
x"ff470",-- -185
x"feee0",-- -274
x"feb70",-- -329
x"fe730",-- -397
x"fe5d0",-- -419
x"febb0",-- -325
x"ff1c0",-- -228
x"ff440",-- -188
x"ff920",-- -110
x"00120",-- 18
x"00730",-- 115
x"00870",-- 135
x"00960",-- 150
x"009d0",-- 157
x"006c0",-- 108
x"00430",-- 67
x"00140",-- 20
x"ffc10",-- -63
x"ff900",-- -112
x"ffc90",-- -55
x"ffd80",-- -40
x"ffb20",-- -78
x"ffbf0",-- -65
x"ffd50",-- -43
x"ffdf0",-- -33
x"ffc10",-- -63
x"ffa30",-- -93
x"ff9e0",-- -98
x"ffb20",-- -78
x"ffb30",-- -77
x"ff680",-- -152
x"ff990",-- -103
x"00070",-- 7
x"000f0",-- 15
x"00140",-- 20
x"00490",-- 73
x"006b0",-- 107
x"00610",-- 97
x"003c0",-- 60
x"00460",-- 70
x"00370",-- 55
x"002b0",-- 43
x"00160",-- 22
x"ffe50",-- -27
x"ffee0",-- -18
x"000c0",-- 12
x"002b0",-- 43
x"002f0",-- 47
x"006b0",-- 107
x"00ad0",-- 173
x"00cb0",-- 203
x"011d0",-- 285
x"013d0",-- 317
x"01350",-- 309
x"01590",-- 345
x"015d0",-- 349
x"01260",-- 294
x"00f20",-- 242
x"00e90",-- 233
x"00bc0",-- 188
x"005f0",-- 95
x"001e0",-- 30
x"ffe50",-- -27
x"ffc90",-- -55
x"ffab0",-- -85
x"ffa90",-- -87
x"ffa90",-- -87
x"ffb80",-- -72
x"ffea0",-- -22
x"fff10",-- -15
x"fffb0",-- -5
x"00230",-- 35
x"00640",-- 100
x"00640",-- 100
x"00300",-- 48
x"00110",-- 17
x"002f0",-- 47
x"002b0",-- 43
x"ffe50",-- -27
x"ffa30",-- -93
x"ffae0",-- -82
x"ffd30",-- -45
x"ffc60",-- -58
x"ffdb0",-- -37
x"ffea0",-- -22
x"ffec0",-- -20
x"ffbd0",-- -67
x"ff630",-- -157
x"ff290",-- -215
x"ff010",-- -255
x"feff0",-- -257
x"fefd0",-- -259
x"fed40",-- -300
x"fedf0",-- -289
x"ff2e0",-- -210
x"ff590",-- -167
x"ff4f0",-- -177
x"ff580",-- -168
x"ffa90",-- -87
x"ffd30",-- -45
x"ffc70",-- -57
x"ffec0",-- -20
x"001c0",-- 28
x"003f0",-- 63
x"002a0",-- 42
x"000c0",-- 12
x"00280",-- 40
x"00410",-- 65
x"00480",-- 72
x"00280",-- 40
x"002b0",-- 43
x"00260",-- 38
x"00030",-- 3
x"ffdb0",-- -37
x"ff970",-- -105
x"ff920",-- -110
x"ff830",-- -125
x"ff710",-- -143
x"ff6a0",-- -150
x"ff6d0",-- -147
x"ff7b0",-- -133
x"ff9e0",-- -98
x"ff9a0",-- -102
x"ff810",-- -127
x"ffae0",-- -82
x"ffdd0",-- -35
x"ffbd0",-- -67
x"ffb70",-- -73
x"ffda0",-- -38
x"fff80",-- -8
x"00050",-- 5
x"00050",-- 5
x"00050",-- 5
x"00320",-- 50
x"00700",-- 112
x"00340",-- 52
x"00000",-- 0
x"00110",-- 17
x"fff80",-- -8
x"ffb80",-- -72
x"ffa60",-- -90
x"ffc60",-- -58
x"ffb30",-- -77
x"ff9e0",-- -98
x"ffa90",-- -87
x"ff970",-- -105
x"ff900",-- -112
x"ff8d0",-- -115
x"ff8d0",-- -115
x"ff940",-- -108
x"ff8d0",-- -115
x"ffa30",-- -93
x"ffd10",-- -47
x"ffe50",-- -27
x"ffce0",-- -50
x"ffdb0",-- -37
x"ffea0",-- -22
x"ffe00",-- -32
x"ffc90",-- -55
x"ffb50",-- -75
x"ffbf0",-- -65
x"ffe40",-- -28
x"fffd0",-- -3
x"00050",-- 5
x"002f0",-- 47
x"00580",-- 88
x"00430",-- 67
x"00160",-- 22
x"00080",-- 8
x"00050",-- 5
x"ffec0",-- -20
x"ffb30",-- -77
x"ff8d0",-- -115
x"ff8b0",-- -117
x"ffa10",-- -95
x"ffb30",-- -77
x"ffc90",-- -55
x"fff40",-- -12
x"001e0",-- 30
x"003c0",-- 60
x"00300",-- 48
x"002f0",-- 47
x"00620",-- 98
x"00660",-- 102
x"00410",-- 65
x"00080",-- 8
x"ffef0",-- -17
x"ffec0",-- -20
x"ffbc0",-- -68
x"ff5d0",-- -163
x"ff470",-- -185
x"ff300",-- -208
x"ff090",-- -247
x"feed0",-- -275
x"ff020",-- -254
x"ff350",-- -203
x"ff1c0",-- -228
x"ff010",-- -255
x"fefa0",-- -262
x"fefd0",-- -259
x"ff1f0",-- -225
x"ff2b0",-- -213
x"ff580",-- -168
x"ffa40",-- -92
x"ffc60",-- -58
x"fff60",-- -10
x"000a0",-- 10
x"00070",-- 7
x"00110",-- 17
x"fffe0",-- -2
x"ffd80",-- -40
x"ffb20",-- -78
x"ff880",-- -120
x"ff880",-- -120
x"ff800",-- -128
x"ff450",-- -187
x"ff100",-- -240
x"ff130",-- -237
x"ff560",-- -170
x"ff650",-- -155
x"ff630",-- -157
x"ff950",-- -107
x"ffcc0",-- -52
x"ffee0",-- -18
x"ffdf0",-- -33
x"ffda0",-- -38
x"00110",-- 17
x"002a0",-- 42
x"ffee0",-- -18
x"ffb20",-- -78
x"ffa80",-- -88
x"ffbc0",-- -68
x"ff860",-- -122
x"ff4a0",-- -182
x"ff540",-- -172
x"ff850",-- -123
x"ff900",-- -112
x"ff7e0",-- -130
x"ff860",-- -122
x"ffae0",-- -82
x"ffcb0",-- -53
x"ffc60",-- -58
x"ffc70",-- -57
x"ffcc0",-- -52
x"fffd0",-- -3
x"00120",-- 18
x"fff80",-- -8
x"fff80",-- -8
x"000c0",-- 12
x"001e0",-- 30
x"000c0",-- 12
x"00140",-- 20
x"001c0",-- 28
x"001b0",-- 27
x"00320",-- 50
x"002f0",-- 47
x"00080",-- 8
x"00110",-- 17
x"00280",-- 40
x"00200",-- 32
x"00000",-- 0
x"00080",-- 8
x"00320",-- 50
x"00200",-- 32
x"00080",-- 8
x"00170",-- 23
x"00490",-- 73
x"00870",-- 135
x"00990",-- 153
x"00a80",-- 168
x"00c60",-- 198
x"00d70",-- 215
x"00c00",-- 192
x"009e0",-- 158
x"00a80",-- 168
x"009b0",-- 155
x"007b0",-- 123
x"00610",-- 97
x"00350",-- 53
x"00370",-- 55
x"00440",-- 68
x"00320",-- 50
x"001c0",-- 28
x"002a0",-- 42
x"00280",-- 40
x"000c0",-- 12
x"001e0",-- 30
x"00440",-- 68
x"00580",-- 88
x"00610",-- 97
x"007a0",-- 122
x"007a0",-- 122
x"00700",-- 112
x"00ac0",-- 172
x"00c30",-- 195
x"00a00",-- 160
x"00940",-- 148
x"008c0",-- 140
x"006e0",-- 110
x"00210",-- 33
x"000c0",-- 12
x"00190",-- 25
x"fffb0",-- -5
x"ffa80",-- -88
x"ff670",-- -153
x"ff7c0",-- -132
x"ff9f0",-- -97
x"ff9f0",-- -97
x"ffb80",-- -72
x"fffe0",-- -2
x"00410",-- 65
x"00440",-- 68
x"006e0",-- 110
x"00c00",-- 192
x"00d20",-- 210
x"00e40",-- 228
x"00d50",-- 213
x"009d0",-- 157
x"007d0",-- 125
x"00840",-- 132
x"00760",-- 118
x"001e0",-- 30
x"ffec0",-- -20
x"ffe50",-- -27
x"ffb70",-- -73
x"ff940",-- -108
x"ff810",-- -127
x"ffa30",-- -93
x"ffa90",-- -87
x"ff6c0",-- -148
x"ff6f0",-- -145
x"ff970",-- -105
x"ffdb0",-- -37
x"00000",-- 0
x"002b0",-- 43
x"00760",-- 118
x"009d0",-- 157
x"00bb0",-- 187
x"00af0",-- 175
x"00a50",-- 165
x"009b0",-- 155
x"00620",-- 98
x"001b0",-- 27
x"fff10",-- -15
x"ffea0",-- -22
x"ffd50",-- -43
x"ffbd0",-- -67
x"ffba0",-- -70
x"ff950",-- -107
x"ff8a0",-- -118
x"ff9e0",-- -98
x"ffba0",-- -70
x"ffad0",-- -83
x"ffc40",-- -60
x"ffe40",-- -28
x"ffdf0",-- -33
x"ffef0",-- -17
x"fffb0",-- -5
x"001e0",-- 30
x"00280",-- 40
x"002d0",-- 45
x"001e0",-- 30
x"00000",-- 0
x"00000",-- 0
x"ffea0",-- -22
x"ffd80",-- -40
x"ffcb0",-- -53
x"ffd60",-- -42
x"fff40",-- -12
x"ffe40",-- -28
x"ffea0",-- -22
x"00000",-- 0
x"000c0",-- 12
x"00050",-- 5
x"000a0",-- 10
x"000f0",-- 15
x"00000",-- 0
x"fffe0",-- -2
x"ffe00",-- -32
x"ffe20",-- -30
x"ffe00",-- -32
x"fffb0",-- -5
x"fff40",-- -12
x"ffd60",-- -42
x"00070",-- 7
x"002a0",-- 42
x"001e0",-- 30
x"000f0",-- 15
x"00190",-- 25
x"00190",-- 25
x"fffb0",-- -5
x"fffb0",-- -5
x"fff90",-- -7
x"00030",-- 3
x"00250",-- 37
x"00370",-- 55
x"00190",-- 25
x"00080",-- 8
x"002b0",-- 43
x"00260",-- 38
x"000f0",-- 15
x"000f0",-- 15
x"00210",-- 33
x"00250",-- 37
x"00000",-- 0
x"00000",-- 0
x"00320",-- 50
x"003a0",-- 58
x"00320",-- 50
x"00200",-- 32
x"00410",-- 65
x"004e0",-- 78
x"002b0",-- 43
x"00280",-- 40
x"002b0",-- 43
x"00120",-- 18
x"ffd80",-- -40
x"ffd30",-- -45
x"ffd80",-- -40
x"ffea0",-- -22
x"ffef0",-- -17
x"00000",-- 0
x"000d0",-- 13
x"00110",-- 17
x"00110",-- 17
x"fffe0",-- -2
x"ffe90",-- -23
x"ffce0",-- -50
x"ffc90",-- -55
x"ffad0",-- -83
x"ff8d0",-- -115
x"ff7e0",-- -130
x"ff9f0",-- -97
x"ffbd0",-- -67
x"ffcb0",-- -53
x"00000",-- 0
x"003f0",-- 63
x"006b0",-- 107
x"007a0",-- 122
x"007d0",-- 125
x"00610",-- 97
x"00520",-- 82
x"00170",-- 23
x"ffd80",-- -40
x"ffb70",-- -73
x"ff9a0",-- -102
x"ff790",-- -135
x"ff830",-- -125
x"ff8d0",-- -115
x"ff920",-- -110
x"ffad0",-- -83
x"ffbc0",-- -68
x"ffd00",-- -48
x"ffdf0",-- -33
x"fff90",-- -7
x"00000",-- 0
x"ffee0",-- -18
x"ffe50",-- -27
x"00030",-- 3
x"00210",-- 33
x"002a0"-- 42
);
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: top PORT MAP (
          clk => clk,
          rstn => rstn,
          i_volume => i_volume,
			 i_agc_enable => i_agc_enable,
          i_SDATA_IN => i_SDATA_IN,
          o_SDATA_out => o_SDATA_out,
          o_SYNC => o_SYNC,
          o_RSTN => o_RSTN,
          i_BIT_CLK => i_BIT_CLK
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 
   i_BIT_CLK_process :process
   begin
		i_BIT_CLK <= '0';
		wait for i_BIT_CLK_period/2;
		i_BIT_CLK <= '1';
		wait for i_BIT_CLK_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin	
		rstn <= '0';
		-- hold reset state for 100 ns.
		wait for 100 ns;	
		rstn <= '1';
		i_volume <= (others => '1');

	wait for i_bit_clk_period*56;
		
		for j in 0 to len-1 loop
			--for k in 0 to 1 loop
				for i in 19 downto 0 loop
					i_sdata_in <= s(j)(i);
					wait for i_bit_clk_period;
				end loop;
				for i in 19 downto 0 loop
					i_sdata_in <= s(j)(i);
					wait for i_bit_clk_period;
				end loop;
			--end loop;
			wait for i_bit_clk_period*216;
		end loop;

		wait;
   end process;

END;
