        when x"12" => gain_n <= x"207"; -- 100dB
        when x"11" => gain_n <= x"28d"; -- 99dB
        when x"10" => gain_n <= x"337"; -- 98dB
        when x"0f" => gain_n <= x"40c"; -- 97dB
        when x"0e" => gain_n <= x"518"; -- 96dB
        when x"0d" => gain_n <= x"66a"; -- 95dB
        when x"0c" => gain_n <= x"813"; -- 94dB
        when x"0b" => gain_n <= x"a2a"; -- 93dB
        when x"0a" => gain_n <= x"ccc"; -- 92dB
        when x"09" => gain_n <= x"101d"; -- 91dB
        when x"08" => gain_n <= x"1449"; -- 90dB
        when x"07" => gain_n <= x"1a1d"; -- 89dB
        when x"06" => gain_n <= x"1d1c"; -- 88dB
        when x"05" => gain_n <= x"2016"; -- 87dB
        when x"04" => gain_n <= x"230d"; -- 86dB
        when x"03" => gain_n <= x"25fe"; -- 85dB
        when x"02" => gain_n <= x"28eb"; -- 84dB
        when x"01" => gain_n <= x"2bd4"; -- 83dB
        when x"00" => gain_n <= x"2eb7"; -- 82dB
        when x"ff" => gain_n <= x"3195"; -- 81dB
        when x"fe" => gain_n <= x"346e"; -- 80dB
        when x"fd" => gain_n <= x"3742"; -- 79dB
        when x"fc" => gain_n <= x"3a10"; -- 78dB
        when x"fb" => gain_n <= x"3cd7"; -- 77dB
        when x"fa" => gain_n <= x"3f99"; -- 76dB
        when x"f9" => gain_n <= x"4254"; -- 75dB
        when x"f8" => gain_n <= x"4508"; -- 74dB
        when x"f7" => gain_n <= x"47b6"; -- 73dB
        when x"f6" => gain_n <= x"4a5c"; -- 72dB
        when x"f5" => gain_n <= x"4cfa"; -- 71dB
        when x"f4" => gain_n <= x"4f91"; -- 70dB
        when x"f3" => gain_n <= x"5220"; -- 69dB
        when x"f2" => gain_n <= x"54a5"; -- 68dB
        when x"f1" => gain_n <= x"5722"; -- 67dB
        when x"f0" => gain_n <= x"5996"; -- 66dB
        when x"ef" => gain_n <= x"5bff"; -- 65dB
        when x"ee" => gain_n <= x"5e5e"; -- 64dB
        when x"ed" => gain_n <= x"60b3"; -- 63dB
        when x"ec" => gain_n <= x"62fc"; -- 62dB
        when x"eb" => gain_n <= x"6539"; -- 61dB
        when x"ea" => gain_n <= x"676a"; -- 60dB
        when x"e9" => gain_n <= x"698e"; -- 59dB
        when x"e8" => gain_n <= x"6ba4"; -- 58dB
        when x"e7" => gain_n <= x"6dab"; -- 57dB
        when x"e6" => gain_n <= x"6fa4"; -- 56dB
        when x"e5" => gain_n <= x"718c"; -- 55dB
        when x"e4" => gain_n <= x"7363"; -- 54dB
        when x"e3" => gain_n <= x"7528"; -- 53dB
        when x"e2" => gain_n <= x"76da"; -- 52dB
        when x"e1" => gain_n <= x"7878"; -- 51dB
        when x"e0" => gain_n <= x"7a01"; -- 50dB
        when x"df" => gain_n <= x"7b73"; -- 49dB
        when x"de" => gain_n <= x"7ccd"; -- 48dB
        when x"dd" => gain_n <= x"7e0d"; -- 47dB
        when x"dc" => gain_n <= x"7f33"; -- 46dB
        when x"db" => gain_n <= x"7fff"; -- 45dB
        when x"da" => gain_n <= x"7fff"; -- 44dB
        when x"d9" => gain_n <= x"7fff"; -- 43dB
        when x"d8" => gain_n <= x"7fff"; -- 42dB
        when x"d7" => gain_n <= x"7fff"; -- 41dB
        when x"d6" => gain_n <= x"7fff"; -- 40dB
        when x"d5" => gain_n <= x"7fff"; -- 39dB
        when x"d4" => gain_n <= x"7fff"; -- 38dB
        when x"d3" => gain_n <= x"7fff"; -- 37dB
        when x"d2" => gain_n <= x"7fff"; -- 36dB
        when x"d1" => gain_n <= x"7fff"; -- 35dB
        when x"d0" => gain_n <= x"7fff"; -- 34dB
        when x"cf" => gain_n <= x"7fff"; -- 33dB
        when x"ce" => gain_n <= x"7fff"; -- 32dB
        when x"cd" => gain_n <= x"7fff"; -- 31dB
        when x"cc" => gain_n <= x"7fff"; -- 30dB
        when x"cb" => gain_n <= x"7fff"; -- 29dB
        when x"ca" => gain_n <= x"7fff"; -- 28dB
        when x"c9" => gain_n <= x"7fff"; -- 27dB
        when x"c8" => gain_n <= x"7fff"; -- 26dB
        when x"c7" => gain_n <= x"7fff"; -- 25dB
        when x"c6" => gain_n <= x"7fff"; -- 24dB
        when x"c5" => gain_n <= x"7fff"; -- 23dB
        when x"c4" => gain_n <= x"7fff"; -- 22dB
        when x"c3" => gain_n <= x"7fff"; -- 21dB
        when x"c2" => gain_n <= x"7fff"; -- 20dB
        when x"c1" => gain_n <= x"7fff"; -- 19dB
        when x"c0" => gain_n <= x"7fff"; -- 18dB
        when x"bf" => gain_n <= x"7fff"; -- 17dB
        when x"be" => gain_n <= x"7fff"; -- 16dB
        when x"bd" => gain_n <= x"7fff"; -- 15dB
        when x"bc" => gain_n <= x"7fff"; -- 14dB
        when x"bb" => gain_n <= x"7fff"; -- 13dB
        when x"ba" => gain_n <= x"7fff"; -- 12dB
        when x"b9" => gain_n <= x"7fff"; -- 11dB
        when x"b8" => gain_n <= x"7fff"; -- 10dB
        when x"b7" => gain_n <= x"7fff"; -- 9dB
        when x"b6" => gain_n <= x"7fff"; -- 8dB
        when x"b5" => gain_n <= x"7fff"; -- 7dB
        when x"b4" => gain_n <= x"7fff"; -- 6dB
        when x"b3" => gain_n <= x"7fff"; -- 5dB
        when x"b2" => gain_n <= x"7fff"; -- 4dB
        when x"b1" => gain_n <= x"7fff"; -- 3dB
        when x"b0" => gain_n <= x"7fff"; -- 2dB
        when x"af" => gain_n <= x"7fff"; -- 1dB
